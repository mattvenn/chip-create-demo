magic
tech sky130A
magscale 1 2
timestamp 1757586453
<< viali >>
rect 24593 47209 24627 47243
rect 5273 47141 5307 47175
rect 22477 47073 22511 47107
rect 5457 47005 5491 47039
rect 5733 47005 5767 47039
rect 22109 47005 22143 47039
rect 10701 45441 10735 45475
rect 10885 45441 10919 45475
rect 10977 45441 11011 45475
rect 11805 45441 11839 45475
rect 11989 45441 12023 45475
rect 13829 45441 13863 45475
rect 13921 45441 13955 45475
rect 14473 45441 14507 45475
rect 14657 45441 14691 45475
rect 16037 45441 16071 45475
rect 17141 45441 17175 45475
rect 17325 45441 17359 45475
rect 19708 45441 19742 45475
rect 17049 45373 17083 45407
rect 18337 45373 18371 45407
rect 19441 45373 19475 45407
rect 20821 45305 20855 45339
rect 10517 45237 10551 45271
rect 11621 45237 11655 45271
rect 13645 45237 13679 45271
rect 14657 45237 14691 45271
rect 14933 45237 14967 45271
rect 15945 45237 15979 45271
rect 17509 45237 17543 45271
rect 17785 45237 17819 45271
rect 10057 45033 10091 45067
rect 16497 45033 16531 45067
rect 19993 45033 20027 45067
rect 10241 44965 10275 44999
rect 11253 44965 11287 44999
rect 15577 44965 15611 44999
rect 10885 44897 10919 44931
rect 13001 44897 13035 44931
rect 15853 44897 15887 44931
rect 7481 44829 7515 44863
rect 8033 44829 8067 44863
rect 8217 44829 8251 44863
rect 10517 44829 10551 44863
rect 10701 44829 10735 44863
rect 10793 44829 10827 44863
rect 11069 44829 11103 44863
rect 11529 44829 11563 44863
rect 14197 44829 14231 44863
rect 17141 44829 17175 44863
rect 19349 44829 19383 44863
rect 9873 44761 9907 44795
rect 10078 44761 10112 44795
rect 12173 44761 12207 44795
rect 14464 44761 14498 44795
rect 17408 44761 17442 44795
rect 6929 44693 6963 44727
rect 7849 44693 7883 44727
rect 8585 44693 8619 44727
rect 12449 44693 12483 44727
rect 18521 44693 18555 44727
rect 9597 44489 9631 44523
rect 11253 44489 11287 44523
rect 14105 44489 14139 44523
rect 14657 44489 14691 44523
rect 20545 44489 20579 44523
rect 6929 44421 6963 44455
rect 7450 44421 7484 44455
rect 10140 44421 10174 44455
rect 15025 44421 15059 44455
rect 4721 44353 4755 44387
rect 4905 44353 4939 44387
rect 6745 44353 6779 44387
rect 9413 44353 9447 44387
rect 9597 44353 9631 44387
rect 12541 44353 12575 44387
rect 12633 44353 12667 44387
rect 12817 44353 12851 44387
rect 13461 44353 13495 44387
rect 14105 44353 14139 44387
rect 14289 44353 14323 44387
rect 16037 44353 16071 44387
rect 16130 44353 16164 44387
rect 16773 44353 16807 44387
rect 17785 44353 17819 44387
rect 18052 44353 18086 44387
rect 20361 44353 20395 44387
rect 20637 44353 20671 44387
rect 6561 44285 6595 44319
rect 7205 44285 7239 44319
rect 9873 44285 9907 44319
rect 11621 44285 11655 44319
rect 11805 44285 11839 44319
rect 11897 44285 11931 44319
rect 11989 44285 12023 44319
rect 12081 44285 12115 44319
rect 13369 44285 13403 44319
rect 15117 44285 15151 44319
rect 15209 44285 15243 44319
rect 17325 44285 17359 44319
rect 19441 44285 19475 44319
rect 13829 44217 13863 44251
rect 16405 44217 16439 44251
rect 19165 44217 19199 44251
rect 20361 44217 20395 44251
rect 4537 44149 4571 44183
rect 8585 44149 8619 44183
rect 13001 44149 13035 44183
rect 20085 44149 20119 44183
rect 21005 44149 21039 44183
rect 7113 43945 7147 43979
rect 9597 43945 9631 43979
rect 12909 43945 12943 43979
rect 13369 43945 13403 43979
rect 18153 43945 18187 43979
rect 20269 43945 20303 43979
rect 20453 43945 20487 43979
rect 13461 43877 13495 43911
rect 17877 43877 17911 43911
rect 9873 43809 9907 43843
rect 12449 43809 12483 43843
rect 13829 43809 13863 43843
rect 14197 43809 14231 43843
rect 14473 43809 14507 43843
rect 15025 43809 15059 43843
rect 20821 43809 20855 43843
rect 4445 43741 4479 43775
rect 8493 43741 8527 43775
rect 9321 43741 9355 43775
rect 9413 43741 9447 43775
rect 11805 43741 11839 43775
rect 11897 43741 11931 43775
rect 11989 43741 12023 43775
rect 12173 43741 12207 43775
rect 12541 43741 12575 43775
rect 12725 43741 12759 43775
rect 14565 43741 14599 43775
rect 16681 43741 16715 43775
rect 16774 43741 16808 43775
rect 17146 43741 17180 43775
rect 17601 43741 17635 43775
rect 17693 43741 17727 43775
rect 18797 43741 18831 43775
rect 19349 43741 19383 43775
rect 19533 43741 19567 43775
rect 19717 43741 19751 43775
rect 19809 43741 19843 43775
rect 20729 43741 20763 43775
rect 20913 43741 20947 43775
rect 4712 43673 4746 43707
rect 8226 43673 8260 43707
rect 10140 43673 10174 43707
rect 11529 43673 11563 43707
rect 15292 43673 15326 43707
rect 16957 43673 16991 43707
rect 17049 43673 17083 43707
rect 17877 43673 17911 43707
rect 20085 43673 20119 43707
rect 5825 43605 5859 43639
rect 11253 43605 11287 43639
rect 16405 43605 16439 43639
rect 17325 43605 17359 43639
rect 20285 43605 20319 43639
rect 21189 43605 21223 43639
rect 11069 43401 11103 43435
rect 13185 43401 13219 43435
rect 15853 43401 15887 43435
rect 16773 43401 16807 43435
rect 20545 43401 20579 43435
rect 10425 43333 10459 43367
rect 13369 43333 13403 43367
rect 6469 43265 6503 43299
rect 10793 43265 10827 43299
rect 10885 43265 10919 43299
rect 11621 43265 11655 43299
rect 12541 43265 12575 43299
rect 13553 43265 13587 43299
rect 14013 43265 14047 43299
rect 16957 43265 16991 43299
rect 17049 43265 17083 43299
rect 17325 43265 17359 43299
rect 17693 43265 17727 43299
rect 17785 43265 17819 43299
rect 18245 43265 18279 43299
rect 18512 43265 18546 43299
rect 14105 43197 14139 43231
rect 15209 43197 15243 43231
rect 19901 43197 19935 43231
rect 14381 43129 14415 43163
rect 17233 43129 17267 43163
rect 19625 43129 19659 43163
rect 7113 43061 7147 43095
rect 12265 43061 12299 43095
rect 12633 43061 12667 43095
rect 17969 43061 18003 43095
rect 11713 42857 11747 42891
rect 12541 42857 12575 42891
rect 16681 42857 16715 42891
rect 18889 42789 18923 42823
rect 10977 42721 11011 42755
rect 12081 42721 12115 42755
rect 14289 42721 14323 42755
rect 14933 42721 14967 42755
rect 15117 42721 15151 42755
rect 18429 42721 18463 42755
rect 18521 42721 18555 42755
rect 19349 42721 19383 42755
rect 19901 42721 19935 42755
rect 5089 42653 5123 42687
rect 11161 42653 11195 42687
rect 11943 42653 11977 42687
rect 12449 42653 12483 42687
rect 12633 42653 12667 42687
rect 14197 42653 14231 42687
rect 14381 42653 14415 42687
rect 14657 42653 14691 42687
rect 15025 42653 15059 42687
rect 16129 42653 16163 42687
rect 16497 42653 16531 42687
rect 18705 42653 18739 42687
rect 5356 42585 5390 42619
rect 11345 42585 11379 42619
rect 16313 42585 16347 42619
rect 16405 42585 16439 42619
rect 6469 42517 6503 42551
rect 14749 42517 14783 42551
rect 15485 42517 15519 42551
rect 17969 42517 18003 42551
rect 5457 42313 5491 42347
rect 19441 42313 19475 42347
rect 5641 42177 5675 42211
rect 5825 42177 5859 42211
rect 6469 42177 6503 42211
rect 19349 42177 19383 42211
rect 19533 42177 19567 42211
rect 7113 41973 7147 42007
rect 19901 41973 19935 42007
rect 6009 41633 6043 41667
rect 5825 41565 5859 41599
rect 13553 41565 13587 41599
rect 5641 41429 5675 41463
rect 13645 41429 13679 41463
rect 7573 41225 7607 41259
rect 7389 41157 7423 41191
rect 4721 41089 4755 41123
rect 4988 41089 5022 41123
rect 7113 41089 7147 41123
rect 7665 41089 7699 41123
rect 7757 41089 7791 41123
rect 6469 41021 6503 41055
rect 6101 40953 6135 40987
rect 7941 40885 7975 40919
rect 6837 40681 6871 40715
rect 8125 40681 8159 40715
rect 9505 40681 9539 40715
rect 16221 40681 16255 40715
rect 8309 40613 8343 40647
rect 6837 40545 6871 40579
rect 7941 40545 7975 40579
rect 6101 40477 6135 40511
rect 6285 40477 6319 40511
rect 6653 40477 6687 40511
rect 6929 40477 6963 40511
rect 8125 40477 8159 40511
rect 10149 40477 10183 40511
rect 16037 40477 16071 40511
rect 7849 40409 7883 40443
rect 15853 40409 15887 40443
rect 5917 40341 5951 40375
rect 7113 40341 7147 40375
rect 7665 40137 7699 40171
rect 9321 40137 9355 40171
rect 10977 40137 11011 40171
rect 11621 40137 11655 40171
rect 16037 40137 16071 40171
rect 7941 40001 7975 40035
rect 8208 40001 8242 40035
rect 9597 40001 9631 40035
rect 9853 40001 9887 40035
rect 11989 40001 12023 40035
rect 14564 40001 14598 40035
rect 14657 40001 14691 40035
rect 15577 40001 15611 40035
rect 7021 39933 7055 39967
rect 11805 39933 11839 39967
rect 11897 39933 11931 39967
rect 12081 39933 12115 39967
rect 18245 39933 18279 39967
rect 15853 39865 15887 39899
rect 14473 39797 14507 39831
rect 16405 39797 16439 39831
rect 18889 39797 18923 39831
rect 7021 39593 7055 39627
rect 7665 39593 7699 39627
rect 9413 39593 9447 39627
rect 16037 39593 16071 39627
rect 10609 39525 10643 39559
rect 15025 39525 15059 39559
rect 5641 39457 5675 39491
rect 7297 39457 7331 39491
rect 8125 39457 8159 39491
rect 9045 39457 9079 39491
rect 9689 39457 9723 39491
rect 11621 39457 11655 39491
rect 12081 39457 12115 39491
rect 15117 39457 15151 39491
rect 18521 39457 18555 39491
rect 5908 39389 5942 39423
rect 7481 39389 7515 39423
rect 9229 39389 9263 39423
rect 10241 39389 10275 39423
rect 10793 39389 10827 39423
rect 10977 39389 11011 39423
rect 11161 39389 11195 39423
rect 11989 39389 12023 39423
rect 15393 39389 15427 39423
rect 15486 39389 15520 39423
rect 15669 39389 15703 39423
rect 15858 39389 15892 39423
rect 16405 39389 16439 39423
rect 18429 39389 18463 39423
rect 18705 39389 18739 39423
rect 18889 39389 18923 39423
rect 19901 39389 19935 39423
rect 10885 39321 10919 39355
rect 14657 39321 14691 39355
rect 15761 39321 15795 39355
rect 8677 39253 8711 39287
rect 17693 39253 17727 39287
rect 19349 39253 19383 39287
rect 7757 39049 7791 39083
rect 8125 39049 8159 39083
rect 13185 39049 13219 39083
rect 17877 39049 17911 39083
rect 20085 39049 20119 39083
rect 7573 38981 7607 39015
rect 8668 38981 8702 39015
rect 20453 38981 20487 39015
rect 7481 38913 7515 38947
rect 7849 38913 7883 38947
rect 8401 38913 8435 38947
rect 10977 38913 11011 38947
rect 13369 38913 13403 38947
rect 13645 38913 13679 38947
rect 13921 38913 13955 38947
rect 14105 38913 14139 38947
rect 15853 38913 15887 38947
rect 15945 38913 15979 38947
rect 16037 38913 16071 38947
rect 16865 38913 16899 38947
rect 19001 38913 19035 38947
rect 19533 38913 19567 38947
rect 19717 38913 19751 38947
rect 19993 38913 20027 38947
rect 20177 38913 20211 38947
rect 20821 38913 20855 38947
rect 7941 38845 7975 38879
rect 10609 38845 10643 38879
rect 11253 38845 11287 38879
rect 12817 38845 12851 38879
rect 14473 38845 14507 38879
rect 15117 38845 15151 38879
rect 19257 38845 19291 38879
rect 9781 38777 9815 38811
rect 11069 38777 11103 38811
rect 13553 38777 13587 38811
rect 10057 38709 10091 38743
rect 11161 38709 11195 38743
rect 12265 38709 12299 38743
rect 14013 38709 14047 38743
rect 15669 38709 15703 38743
rect 19533 38709 19567 38743
rect 9045 38505 9079 38539
rect 9689 38505 9723 38539
rect 17141 38505 17175 38539
rect 17325 38505 17359 38539
rect 11069 38437 11103 38471
rect 15577 38437 15611 38471
rect 18981 38437 19015 38471
rect 9413 38369 9447 38403
rect 12449 38369 12483 38403
rect 14197 38369 14231 38403
rect 17601 38369 17635 38403
rect 19349 38369 19383 38403
rect 1501 38301 1535 38335
rect 1961 38301 1995 38335
rect 9229 38301 9263 38335
rect 10517 38301 10551 38335
rect 10793 38301 10827 38335
rect 12182 38301 12216 38335
rect 12817 38301 12851 38335
rect 13001 38301 13035 38335
rect 13093 38301 13127 38335
rect 13185 38301 13219 38335
rect 15853 38301 15887 38335
rect 16037 38301 16071 38335
rect 10701 38233 10735 38267
rect 13461 38233 13495 38267
rect 14442 38233 14476 38267
rect 16497 38233 16531 38267
rect 16957 38233 16991 38267
rect 17173 38233 17207 38267
rect 17868 38233 17902 38267
rect 1685 38165 1719 38199
rect 10333 38165 10367 38199
rect 15945 38165 15979 38199
rect 19993 38165 20027 38199
rect 10885 37961 10919 37995
rect 12265 37961 12299 37995
rect 13461 37961 13495 37995
rect 15025 37961 15059 37995
rect 16405 37961 16439 37995
rect 18613 37961 18647 37995
rect 19533 37961 19567 37995
rect 9198 37893 9232 37927
rect 13737 37893 13771 37927
rect 14381 37893 14415 37927
rect 15301 37893 15335 37927
rect 15393 37893 15427 37927
rect 16129 37893 16163 37927
rect 2697 37825 2731 37859
rect 3157 37825 3191 37859
rect 3413 37825 3447 37859
rect 8677 37825 8711 37859
rect 11069 37825 11103 37859
rect 11253 37825 11287 37859
rect 11621 37825 11655 37859
rect 11805 37825 11839 37859
rect 11897 37825 11931 37859
rect 11989 37825 12023 37859
rect 14197 37825 14231 37859
rect 14473 37825 14507 37859
rect 14565 37825 14599 37859
rect 15204 37825 15238 37859
rect 15576 37825 15610 37859
rect 15669 37825 15703 37859
rect 16405 37825 16439 37859
rect 18245 37825 18279 37859
rect 19717 37825 19751 37859
rect 2513 37757 2547 37791
rect 2881 37757 2915 37791
rect 5089 37757 5123 37791
rect 8953 37757 8987 37791
rect 12817 37757 12851 37791
rect 17325 37757 17359 37791
rect 19165 37757 19199 37791
rect 19901 37757 19935 37791
rect 4537 37689 4571 37723
rect 7389 37689 7423 37723
rect 14749 37689 14783 37723
rect 16313 37689 16347 37723
rect 16773 37689 16807 37723
rect 5641 37621 5675 37655
rect 10333 37621 10367 37655
rect 17693 37621 17727 37655
rect 12633 37417 12667 37451
rect 13737 37417 13771 37451
rect 14473 37417 14507 37451
rect 18061 37417 18095 37451
rect 18429 37417 18463 37451
rect 16221 37349 16255 37383
rect 9045 37281 9079 37315
rect 10885 37281 10919 37315
rect 11621 37281 11655 37315
rect 12265 37281 12299 37315
rect 12817 37281 12851 37315
rect 14933 37281 14967 37315
rect 17601 37281 17635 37315
rect 17969 37281 18003 37315
rect 4997 37213 5031 37247
rect 7021 37213 7055 37247
rect 10977 37213 11011 37247
rect 12909 37213 12943 37247
rect 13553 37213 13587 37247
rect 14657 37213 14691 37247
rect 14749 37213 14783 37247
rect 15025 37213 15059 37247
rect 15393 37213 15427 37247
rect 17345 37213 17379 37247
rect 18245 37213 18279 37247
rect 5264 37145 5298 37179
rect 15945 37145 15979 37179
rect 6377 37077 6411 37111
rect 11345 37077 11379 37111
rect 5089 36873 5123 36907
rect 12909 36873 12943 36907
rect 16973 36873 17007 36907
rect 17141 36873 17175 36907
rect 15761 36805 15795 36839
rect 16773 36805 16807 36839
rect 5273 36737 5307 36771
rect 5457 36737 5491 36771
rect 12265 36737 12299 36771
rect 12449 36737 12483 36771
rect 13001 36737 13035 36771
rect 15669 36737 15703 36771
rect 15945 36737 15979 36771
rect 7021 36669 7055 36703
rect 12449 36601 12483 36635
rect 15945 36601 15979 36635
rect 6469 36533 6503 36567
rect 16957 36533 16991 36567
rect 5273 36125 5307 36159
rect 7481 36125 7515 36159
rect 5540 36057 5574 36091
rect 4905 35989 4939 36023
rect 6653 35989 6687 36023
rect 6929 35989 6963 36023
rect 4537 35785 4571 35819
rect 6469 35785 6503 35819
rect 16221 35785 16255 35819
rect 16773 35785 16807 35819
rect 16037 35717 16071 35751
rect 3893 35649 3927 35683
rect 4353 35649 4387 35683
rect 4905 35649 4939 35683
rect 4997 35649 5031 35683
rect 7582 35649 7616 35683
rect 7849 35649 7883 35683
rect 16313 35649 16347 35683
rect 4169 35581 4203 35615
rect 6101 35581 6135 35615
rect 5181 35513 5215 35547
rect 5457 35445 5491 35479
rect 16037 35445 16071 35479
rect 5365 35241 5399 35275
rect 11713 35241 11747 35275
rect 16957 35241 16991 35275
rect 14841 35173 14875 35207
rect 18061 35173 18095 35207
rect 5273 35105 5307 35139
rect 6653 35105 6687 35139
rect 9689 35105 9723 35139
rect 5089 35037 5123 35071
rect 5641 35037 5675 35071
rect 6009 35037 6043 35071
rect 6469 35037 6503 35071
rect 6745 35037 6779 35071
rect 7113 35037 7147 35071
rect 9229 35037 9263 35071
rect 9413 35037 9447 35071
rect 11897 35037 11931 35071
rect 12173 35037 12207 35071
rect 16589 35037 16623 35071
rect 5365 34969 5399 35003
rect 5825 34969 5859 35003
rect 5917 34969 5951 35003
rect 9045 34969 9079 35003
rect 4905 34901 4939 34935
rect 6193 34901 6227 34935
rect 6837 34901 6871 34935
rect 7021 34901 7055 34935
rect 12081 34901 12115 34935
rect 16037 34901 16071 34935
rect 7021 34697 7055 34731
rect 13001 34697 13035 34731
rect 14289 34697 14323 34731
rect 16221 34697 16255 34731
rect 10517 34629 10551 34663
rect 12081 34629 12115 34663
rect 12633 34629 12667 34663
rect 16773 34629 16807 34663
rect 5089 34561 5123 34595
rect 5273 34561 5307 34595
rect 6653 34561 6687 34595
rect 6745 34561 6779 34595
rect 6837 34561 6871 34595
rect 7297 34561 7331 34595
rect 8861 34561 8895 34595
rect 9873 34561 9907 34595
rect 10057 34561 10091 34595
rect 10701 34561 10735 34595
rect 12265 34561 12299 34595
rect 14197 34561 14231 34595
rect 14841 34561 14875 34595
rect 14933 34561 14967 34595
rect 15117 34561 15151 34595
rect 15577 34561 15611 34595
rect 5549 34493 5583 34527
rect 6469 34493 6503 34527
rect 9413 34493 9447 34527
rect 9781 34493 9815 34527
rect 9965 34493 9999 34527
rect 10241 34493 10275 34527
rect 10885 34493 10919 34527
rect 19441 34493 19475 34527
rect 4905 34357 4939 34391
rect 7941 34357 7975 34391
rect 15301 34357 15335 34391
rect 18061 34357 18095 34391
rect 18797 34357 18831 34391
rect 5641 34153 5675 34187
rect 6377 34153 6411 34187
rect 8677 34153 8711 34187
rect 10425 34153 10459 34187
rect 16313 34153 16347 34187
rect 17785 34153 17819 34187
rect 10977 34085 11011 34119
rect 13185 34017 13219 34051
rect 17877 34017 17911 34051
rect 4261 33949 4295 33983
rect 6929 33949 6963 33983
rect 7297 33949 7331 33983
rect 9045 33949 9079 33983
rect 9301 33949 9335 33983
rect 10701 33949 10735 33983
rect 11253 33949 11287 33983
rect 11529 33949 11563 33983
rect 12541 33949 12575 33983
rect 12633 33949 12667 33983
rect 12725 33949 12759 33983
rect 12909 33949 12943 33983
rect 14473 33949 14507 33983
rect 14657 33949 14691 33983
rect 14933 33949 14967 33983
rect 16773 33949 16807 33983
rect 17969 33949 18003 33983
rect 18797 33949 18831 33983
rect 19349 33949 19383 33983
rect 22201 33949 22235 33983
rect 25053 33949 25087 33983
rect 4528 33881 4562 33915
rect 7564 33881 7598 33915
rect 15200 33881 15234 33915
rect 17509 33881 17543 33915
rect 17601 33881 17635 33915
rect 12265 33813 12299 33847
rect 13829 33813 13863 33847
rect 14565 33813 14599 33847
rect 18245 33813 18279 33847
rect 19993 33813 20027 33847
rect 21649 33813 21683 33847
rect 24501 33813 24535 33847
rect 9137 33609 9171 33643
rect 10057 33609 10091 33643
rect 11253 33609 11287 33643
rect 16405 33609 16439 33643
rect 19165 33609 19199 33643
rect 19533 33609 19567 33643
rect 7113 33541 7147 33575
rect 10174 33541 10208 33575
rect 11713 33541 11747 33575
rect 15270 33541 15304 33575
rect 24400 33541 24434 33575
rect 6009 33473 6043 33507
rect 9689 33473 9723 33507
rect 9965 33473 9999 33507
rect 12449 33473 12483 33507
rect 14013 33473 14047 33507
rect 14473 33473 14507 33507
rect 15025 33473 15059 33507
rect 17785 33473 17819 33507
rect 18052 33473 18086 33507
rect 19441 33473 19475 33507
rect 19625 33473 19659 33507
rect 21097 33473 21131 33507
rect 21373 33473 21407 33507
rect 21557 33473 21591 33507
rect 21925 33473 21959 33507
rect 22181 33473 22215 33507
rect 23765 33473 23799 33507
rect 10609 33405 10643 33439
rect 14749 33405 14783 33439
rect 21465 33405 21499 33439
rect 24133 33405 24167 33439
rect 26341 33405 26375 33439
rect 12081 33337 12115 33371
rect 13369 33337 13403 33371
rect 14657 33337 14691 33371
rect 25513 33337 25547 33371
rect 5457 33269 5491 33303
rect 8401 33269 8435 33303
rect 10333 33269 10367 33303
rect 12173 33269 12207 33303
rect 13093 33269 13127 33303
rect 14289 33269 14323 33303
rect 23305 33269 23339 33303
rect 23673 33269 23707 33303
rect 25789 33269 25823 33303
rect 5733 33065 5767 33099
rect 5917 33065 5951 33099
rect 10885 33065 10919 33099
rect 12449 33065 12483 33099
rect 14473 33065 14507 33099
rect 16313 33065 16347 33099
rect 17509 33065 17543 33099
rect 19441 33065 19475 33099
rect 21741 33065 21775 33099
rect 23765 33065 23799 33099
rect 6193 32997 6227 33031
rect 9597 32997 9631 33031
rect 15945 32997 15979 33031
rect 17877 32997 17911 33031
rect 18245 32997 18279 33031
rect 5549 32929 5583 32963
rect 9321 32929 9355 32963
rect 10241 32929 10275 32963
rect 11897 32929 11931 32963
rect 13829 32929 13863 32963
rect 18705 32929 18739 32963
rect 21189 32929 21223 32963
rect 21465 32929 21499 32963
rect 22201 32929 22235 32963
rect 22293 32929 22327 32963
rect 23213 32929 23247 32963
rect 25697 32929 25731 32963
rect 5457 32861 5491 32895
rect 5733 32861 5767 32895
rect 6745 32861 6779 32895
rect 9229 32861 9263 32895
rect 11805 32861 11839 32895
rect 13573 32861 13607 32895
rect 14197 32861 14231 32895
rect 14289 32861 14323 32895
rect 15669 32861 15703 32895
rect 17693 32861 17727 32895
rect 17969 32861 18003 32895
rect 18613 32861 18647 32895
rect 19349 32861 19383 32895
rect 19533 32861 19567 32895
rect 19993 32861 20027 32895
rect 21097 32861 21131 32895
rect 22109 32861 22143 32895
rect 25145 32861 25179 32895
rect 25789 32861 25823 32895
rect 7113 32793 7147 32827
rect 14473 32793 14507 32827
rect 14841 32793 14875 32827
rect 15945 32793 15979 32827
rect 12173 32725 12207 32759
rect 15761 32725 15795 32759
rect 19901 32725 19935 32759
rect 24501 32725 24535 32759
rect 25421 32725 25455 32759
rect 6469 32521 6503 32555
rect 10057 32521 10091 32555
rect 11253 32521 11287 32555
rect 11989 32521 12023 32555
rect 17417 32521 17451 32555
rect 21925 32521 21959 32555
rect 23857 32521 23891 32555
rect 24225 32521 24259 32555
rect 25145 32521 25179 32555
rect 5273 32453 5307 32487
rect 23949 32453 23983 32487
rect 5549 32385 5583 32419
rect 5753 32385 5787 32419
rect 7593 32385 7627 32419
rect 9873 32385 9907 32419
rect 10057 32385 10091 32419
rect 10885 32385 10919 32419
rect 11069 32385 11103 32419
rect 11621 32385 11655 32419
rect 11805 32385 11839 32419
rect 12449 32385 12483 32419
rect 12716 32385 12750 32419
rect 15025 32385 15059 32419
rect 15292 32385 15326 32419
rect 18889 32385 18923 32419
rect 19165 32385 19199 32419
rect 22293 32385 22327 32419
rect 22937 32385 22971 32419
rect 23213 32385 23247 32419
rect 23673 32385 23707 32419
rect 24593 32385 24627 32419
rect 25053 32385 25087 32419
rect 25237 32385 25271 32419
rect 25697 32385 25731 32419
rect 27077 32385 27111 32419
rect 7849 32317 7883 32351
rect 10793 32317 10827 32351
rect 16773 32317 16807 32351
rect 22201 32317 22235 32351
rect 23581 32317 23615 32351
rect 24685 32317 24719 32351
rect 28273 32317 28307 32351
rect 13829 32249 13863 32283
rect 16405 32249 16439 32283
rect 18705 32249 18739 32283
rect 1501 32181 1535 32215
rect 5917 32181 5951 32215
rect 11805 32181 11839 32215
rect 19073 32181 19107 32215
rect 22753 32181 22787 32215
rect 23121 32181 23155 32215
rect 23581 32181 23615 32215
rect 25605 32181 25639 32215
rect 7021 31977 7055 32011
rect 7941 31977 7975 32011
rect 12725 31977 12759 32011
rect 15393 31977 15427 32011
rect 16681 31977 16715 32011
rect 18613 31977 18647 32011
rect 19901 31977 19935 32011
rect 21189 31977 21223 32011
rect 22293 31977 22327 32011
rect 6745 31909 6779 31943
rect 7573 31841 7607 31875
rect 8585 31841 8619 31875
rect 16773 31841 16807 31875
rect 19533 31841 19567 31875
rect 19717 31841 19751 31875
rect 20637 31841 20671 31875
rect 21005 31841 21039 31875
rect 21833 31841 21867 31875
rect 22937 31841 22971 31875
rect 5365 31773 5399 31807
rect 8125 31773 8159 31807
rect 8309 31773 8343 31807
rect 12633 31773 12667 31807
rect 12817 31773 12851 31807
rect 16037 31773 16071 31807
rect 16313 31773 16347 31807
rect 16497 31773 16531 31807
rect 18797 31773 18831 31807
rect 18889 31773 18923 31807
rect 19441 31773 19475 31807
rect 19625 31773 19659 31807
rect 20545 31773 20579 31807
rect 20729 31773 20763 31807
rect 21465 31773 21499 31807
rect 21925 31773 21959 31807
rect 22017 31773 22051 31807
rect 22109 31773 22143 31807
rect 22569 31773 22603 31807
rect 22753 31773 22787 31807
rect 24133 31773 24167 31807
rect 28457 31773 28491 31807
rect 5632 31705 5666 31739
rect 18613 31705 18647 31739
rect 21373 31705 21407 31739
rect 7849 31433 7883 31467
rect 22293 31433 22327 31467
rect 21925 31365 21959 31399
rect 22109 31365 22143 31399
rect 6469 31297 6503 31331
rect 6653 31297 6687 31331
rect 7205 31297 7239 31331
rect 21189 31297 21223 31331
rect 21281 31229 21315 31263
rect 21557 31161 21591 31195
rect 6837 31093 6871 31127
rect 5549 30889 5583 30923
rect 18613 30889 18647 30923
rect 6673 30685 6707 30719
rect 6929 30685 6963 30719
rect 18797 30685 18831 30719
rect 18889 30685 18923 30719
rect 7297 30549 7331 30583
rect 17601 30549 17635 30583
rect 17877 30277 17911 30311
rect 18245 30277 18279 30311
rect 18429 30277 18463 30311
rect 24225 30277 24259 30311
rect 1501 30209 1535 30243
rect 1961 30209 1995 30243
rect 17325 30209 17359 30243
rect 17509 30209 17543 30243
rect 17785 30209 17819 30243
rect 17969 30209 18003 30243
rect 23765 30209 23799 30243
rect 23857 30209 23891 30243
rect 24041 30209 24075 30243
rect 9965 30141 9999 30175
rect 18889 30141 18923 30175
rect 19441 30141 19475 30175
rect 1685 30005 1719 30039
rect 8769 30005 8803 30039
rect 9413 30005 9447 30039
rect 17509 30005 17543 30039
rect 18613 30005 18647 30039
rect 10701 29801 10735 29835
rect 15485 29801 15519 29835
rect 18981 29801 19015 29835
rect 19349 29801 19383 29835
rect 24593 29801 24627 29835
rect 9045 29733 9079 29767
rect 8309 29665 8343 29699
rect 11253 29665 11287 29699
rect 17601 29665 17635 29699
rect 19809 29665 19843 29699
rect 19901 29665 19935 29699
rect 1501 29597 1535 29631
rect 8493 29597 8527 29631
rect 10425 29597 10459 29631
rect 17857 29597 17891 29631
rect 23857 29597 23891 29631
rect 23949 29597 23983 29631
rect 8677 29529 8711 29563
rect 10158 29529 10192 29563
rect 19717 29461 19751 29495
rect 24133 29461 24167 29495
rect 9873 29257 9907 29291
rect 18337 29257 18371 29291
rect 26709 29257 26743 29291
rect 10986 29189 11020 29223
rect 12633 29189 12667 29223
rect 14381 29189 14415 29223
rect 22937 29189 22971 29223
rect 23121 29189 23155 29223
rect 24869 29189 24903 29223
rect 3801 29121 3835 29155
rect 7665 29121 7699 29155
rect 8125 29121 8159 29155
rect 9137 29121 9171 29155
rect 13001 29121 13035 29155
rect 13277 29121 13311 29155
rect 13737 29121 13771 29155
rect 13921 29121 13955 29155
rect 14197 29121 14231 29155
rect 15117 29121 15151 29155
rect 15301 29121 15335 29155
rect 15853 29121 15887 29155
rect 16773 29121 16807 29155
rect 16957 29121 16991 29155
rect 18705 29121 18739 29155
rect 19165 29121 19199 29155
rect 23765 29121 23799 29155
rect 25329 29121 25363 29155
rect 25596 29121 25630 29155
rect 3617 29053 3651 29087
rect 4353 29053 4387 29087
rect 7941 29053 7975 29087
rect 8585 29053 8619 29087
rect 11253 29053 11287 29087
rect 12173 29053 12207 29087
rect 15209 29053 15243 29087
rect 15945 29053 15979 29087
rect 16865 29053 16899 29087
rect 18613 29053 18647 29087
rect 23673 29053 23707 29087
rect 24409 29053 24443 29087
rect 3985 28985 4019 29019
rect 8309 28985 8343 29019
rect 13829 28985 13863 29019
rect 14565 28985 14599 29019
rect 16221 28985 16255 29019
rect 23305 28985 23339 29019
rect 24501 28985 24535 29019
rect 11621 28917 11655 28951
rect 19809 28917 19843 28951
rect 24041 28917 24075 28951
rect 8677 28713 8711 28747
rect 11253 28713 11287 28747
rect 11621 28713 11655 28747
rect 15945 28713 15979 28747
rect 17785 28713 17819 28747
rect 26065 28713 26099 28747
rect 5917 28645 5951 28679
rect 17693 28645 17727 28679
rect 21189 28645 21223 28679
rect 6377 28577 6411 28611
rect 7941 28577 7975 28611
rect 9873 28577 9907 28611
rect 15209 28577 15243 28611
rect 17325 28577 17359 28611
rect 17601 28577 17635 28611
rect 20361 28577 20395 28611
rect 21649 28577 21683 28611
rect 21741 28577 21775 28611
rect 25421 28577 25455 28611
rect 4537 28509 4571 28543
rect 7757 28509 7791 28543
rect 8401 28509 8435 28543
rect 8493 28509 8527 28543
rect 10140 28509 10174 28543
rect 12081 28509 12115 28543
rect 14197 28509 14231 28543
rect 14473 28509 14507 28543
rect 14657 28509 14691 28543
rect 16589 28509 16623 28543
rect 16865 28509 16899 28543
rect 17141 28509 17175 28543
rect 17877 28509 17911 28543
rect 19533 28509 19567 28543
rect 23305 28509 23339 28543
rect 23581 28509 23615 28543
rect 25053 28509 25087 28543
rect 4804 28441 4838 28475
rect 7297 28441 7331 28475
rect 8677 28441 8711 28475
rect 9045 28441 9079 28475
rect 9229 28441 9263 28475
rect 12348 28441 12382 28475
rect 14933 28441 14967 28475
rect 16957 28441 16991 28475
rect 23857 28441 23891 28475
rect 6929 28373 6963 28407
rect 7573 28373 7607 28407
rect 8217 28373 8251 28407
rect 9321 28373 9355 28407
rect 9413 28373 9447 28407
rect 9597 28373 9631 28407
rect 13461 28373 13495 28407
rect 19441 28373 19475 28407
rect 20913 28373 20947 28407
rect 21557 28373 21591 28407
rect 24501 28373 24535 28407
rect 10057 28169 10091 28203
rect 10241 28169 10275 28203
rect 10885 28169 10919 28203
rect 13001 28169 13035 28203
rect 15393 28169 15427 28203
rect 16129 28169 16163 28203
rect 17785 28169 17819 28203
rect 22109 28169 22143 28203
rect 24041 28169 24075 28203
rect 24501 28169 24535 28203
rect 25237 28169 25271 28203
rect 14105 28101 14139 28135
rect 6101 28033 6135 28067
rect 6653 28033 6687 28067
rect 6837 28033 6871 28067
rect 7472 28033 7506 28067
rect 9965 28033 9999 28067
rect 10333 28033 10367 28067
rect 11069 28033 11103 28067
rect 11621 28033 11655 28067
rect 11888 28033 11922 28067
rect 13461 28033 13495 28067
rect 16773 28033 16807 28067
rect 17141 28033 17175 28067
rect 17509 28033 17543 28067
rect 17969 28033 18003 28067
rect 20913 28033 20947 28067
rect 21097 28033 21131 28067
rect 21373 28033 21407 28067
rect 22753 28033 22787 28067
rect 23305 28033 23339 28067
rect 23489 28033 23523 28067
rect 24133 28033 24167 28067
rect 24869 28033 24903 28067
rect 24961 28033 24995 28067
rect 7205 27965 7239 27999
rect 9413 27965 9447 27999
rect 10425 27965 10459 27999
rect 11253 27965 11287 27999
rect 13369 27965 13403 27999
rect 18153 27965 18187 27999
rect 20637 27965 20671 27999
rect 23857 27965 23891 27999
rect 8585 27897 8619 27931
rect 13829 27897 13863 27931
rect 6469 27829 6503 27863
rect 8861 27829 8895 27863
rect 10609 27829 10643 27863
rect 20913 27829 20947 27863
rect 21465 27829 21499 27863
rect 23489 27829 23523 27863
rect 8493 27625 8527 27659
rect 9413 27625 9447 27659
rect 12173 27625 12207 27659
rect 12725 27625 12759 27659
rect 14197 27625 14231 27659
rect 17693 27625 17727 27659
rect 22201 27625 22235 27659
rect 25145 27625 25179 27659
rect 7849 27557 7883 27591
rect 8677 27557 8711 27591
rect 16497 27557 16531 27591
rect 17509 27557 17543 27591
rect 24133 27557 24167 27591
rect 8401 27489 8435 27523
rect 10333 27489 10367 27523
rect 13277 27489 13311 27523
rect 14841 27489 14875 27523
rect 16957 27489 16991 27523
rect 17049 27489 17083 27523
rect 24501 27489 24535 27523
rect 6469 27421 6503 27455
rect 8217 27421 8251 27455
rect 8493 27421 8527 27455
rect 10057 27421 10091 27455
rect 11529 27421 11563 27455
rect 16865 27421 16899 27455
rect 18153 27421 18187 27455
rect 20821 27421 20855 27455
rect 22753 27421 22787 27455
rect 23020 27421 23054 27455
rect 28457 27421 28491 27455
rect 6736 27353 6770 27387
rect 15108 27353 15142 27387
rect 17661 27353 17695 27387
rect 17877 27353 17911 27387
rect 21066 27353 21100 27387
rect 10977 27285 11011 27319
rect 16221 27285 16255 27319
rect 18245 27285 18279 27319
rect 8401 27081 8435 27115
rect 10057 27081 10091 27115
rect 11069 27081 11103 27115
rect 12081 27081 12115 27115
rect 12817 27081 12851 27115
rect 13461 27081 13495 27115
rect 17417 27081 17451 27115
rect 25145 27081 25179 27115
rect 10701 27013 10735 27047
rect 10793 27013 10827 27047
rect 22201 27013 22235 27047
rect 22293 27013 22327 27047
rect 23121 27013 23155 27047
rect 7021 26945 7055 26979
rect 7288 26945 7322 26979
rect 8677 26945 8711 26979
rect 8944 26945 8978 26979
rect 10517 26945 10551 26979
rect 10885 26945 10919 26979
rect 12265 26945 12299 26979
rect 12449 26945 12483 26979
rect 13277 26945 13311 26979
rect 13645 26945 13679 26979
rect 13829 26945 13863 26979
rect 14197 26945 14231 26979
rect 14749 26945 14783 26979
rect 16405 26945 16439 26979
rect 16773 26945 16807 26979
rect 18337 26945 18371 26979
rect 18429 26945 18463 26979
rect 18613 26945 18647 26979
rect 21925 26945 21959 26979
rect 22018 26945 22052 26979
rect 22390 26945 22424 26979
rect 22845 26945 22879 26979
rect 23029 26945 23063 26979
rect 23213 26945 23247 26979
rect 23765 26945 23799 26979
rect 23949 26945 23983 26979
rect 24041 26945 24075 26979
rect 24317 26945 24351 26979
rect 25237 26945 25271 26979
rect 15025 26877 15059 26911
rect 16313 26877 16347 26911
rect 24133 26877 24167 26911
rect 24501 26877 24535 26911
rect 24869 26877 24903 26911
rect 14473 26809 14507 26843
rect 22569 26809 22603 26843
rect 23397 26809 23431 26843
rect 13645 26741 13679 26775
rect 18797 26741 18831 26775
rect 24869 26741 24903 26775
rect 24961 26741 24995 26775
rect 8125 26537 8159 26571
rect 13829 26537 13863 26571
rect 17693 26537 17727 26571
rect 17969 26537 18003 26571
rect 20637 26537 20671 26571
rect 22661 26537 22695 26571
rect 8493 26401 8527 26435
rect 9597 26401 9631 26435
rect 18429 26401 18463 26435
rect 20177 26401 20211 26435
rect 20269 26401 20303 26435
rect 8309 26333 8343 26367
rect 12449 26333 12483 26367
rect 17141 26333 17175 26367
rect 17233 26333 17267 26367
rect 17417 26333 17451 26367
rect 17509 26333 17543 26367
rect 18153 26333 18187 26367
rect 18245 26333 18279 26367
rect 18521 26333 18555 26367
rect 19901 26333 19935 26367
rect 20085 26333 20119 26367
rect 20453 26333 20487 26367
rect 22477 26333 22511 26367
rect 12716 26265 12750 26299
rect 22293 26265 22327 26299
rect 9045 26197 9079 26231
rect 9045 25993 9079 26027
rect 12725 25993 12759 26027
rect 13369 25993 13403 26027
rect 18797 25993 18831 26027
rect 19073 25925 19107 25959
rect 9229 25857 9263 25891
rect 9321 25857 9355 25891
rect 12909 25857 12943 25891
rect 13093 25857 13127 25891
rect 18981 25857 19015 25891
rect 19165 25857 19199 25891
rect 19349 25857 19383 25891
rect 13921 25789 13955 25823
rect 25789 25789 25823 25823
rect 8677 25653 8711 25687
rect 9781 25653 9815 25687
rect 12449 25653 12483 25687
rect 25237 25653 25271 25687
rect 21097 25449 21131 25483
rect 19809 25245 19843 25279
rect 19993 25245 20027 25279
rect 20913 25177 20947 25211
rect 19901 25109 19935 25143
rect 21113 25109 21147 25143
rect 21281 25109 21315 25143
rect 18261 24905 18295 24939
rect 18061 24837 18095 24871
rect 21557 24837 21591 24871
rect 23397 24837 23431 24871
rect 23597 24837 23631 24871
rect 12173 24769 12207 24803
rect 12440 24769 12474 24803
rect 19533 24769 19567 24803
rect 20453 24769 20487 24803
rect 22109 24769 22143 24803
rect 22845 24769 22879 24803
rect 23121 24769 23155 24803
rect 19809 24701 19843 24735
rect 20177 24701 20211 24735
rect 21005 24701 21039 24735
rect 22385 24701 22419 24735
rect 13553 24633 13587 24667
rect 18429 24633 18463 24667
rect 19717 24633 19751 24667
rect 22293 24633 22327 24667
rect 18245 24565 18279 24599
rect 19349 24565 19383 24599
rect 20269 24565 20303 24599
rect 20637 24565 20671 24599
rect 21925 24565 21959 24599
rect 22661 24565 22695 24599
rect 23029 24565 23063 24599
rect 23581 24565 23615 24599
rect 23765 24565 23799 24599
rect 11989 24361 12023 24395
rect 21465 24361 21499 24395
rect 24777 24293 24811 24327
rect 17049 24225 17083 24259
rect 18245 24225 18279 24259
rect 20637 24225 20671 24259
rect 23213 24225 23247 24259
rect 23949 24225 23983 24259
rect 1501 24157 1535 24191
rect 11069 24157 11103 24191
rect 12633 24157 12667 24191
rect 17509 24157 17543 24191
rect 17693 24157 17727 24191
rect 17785 24157 17819 24191
rect 18797 24157 18831 24191
rect 19349 24157 19383 24191
rect 22109 24157 22143 24191
rect 23765 24157 23799 24191
rect 24501 24157 24535 24191
rect 24777 24089 24811 24123
rect 25053 24089 25087 24123
rect 10425 24021 10459 24055
rect 16405 24021 16439 24055
rect 17325 24021 17359 24055
rect 19993 24021 20027 24055
rect 21189 24021 21223 24055
rect 22661 24021 22695 24055
rect 23581 24021 23615 24055
rect 24593 24021 24627 24055
rect 10057 23817 10091 23851
rect 12265 23817 12299 23851
rect 16227 23817 16261 23851
rect 18153 23817 18187 23851
rect 20085 23817 20119 23851
rect 23489 23817 23523 23851
rect 25237 23817 25271 23851
rect 16313 23749 16347 23783
rect 17040 23749 17074 23783
rect 19542 23749 19576 23783
rect 8933 23681 8967 23715
rect 10517 23681 10551 23715
rect 10609 23681 10643 23715
rect 12449 23681 12483 23715
rect 12541 23681 12575 23715
rect 13461 23681 13495 23715
rect 13921 23681 13955 23715
rect 15669 23681 15703 23715
rect 15853 23681 15887 23715
rect 16129 23681 16163 23715
rect 16405 23681 16439 23715
rect 19809 23681 19843 23715
rect 21198 23681 21232 23715
rect 21465 23681 21499 23715
rect 23857 23681 23891 23715
rect 24124 23681 24158 23715
rect 8677 23613 8711 23647
rect 12081 23613 12115 23647
rect 12173 23613 12207 23647
rect 13277 23613 13311 23647
rect 16773 23613 16807 23647
rect 22477 23613 22511 23647
rect 22845 23613 22879 23647
rect 1501 23477 1535 23511
rect 10333 23477 10367 23511
rect 10977 23477 11011 23511
rect 12725 23477 12759 23511
rect 13645 23477 13679 23511
rect 15669 23477 15703 23511
rect 18429 23477 18463 23511
rect 21925 23477 21959 23511
rect 11989 23273 12023 23307
rect 13737 23273 13771 23307
rect 20729 23273 20763 23307
rect 21189 23273 21223 23307
rect 22845 23273 22879 23307
rect 23489 23273 23523 23307
rect 24501 23273 24535 23307
rect 24869 23273 24903 23307
rect 12449 23205 12483 23239
rect 12541 23205 12575 23239
rect 14289 23205 14323 23239
rect 16957 23205 16991 23239
rect 17969 23205 18003 23239
rect 15577 23137 15611 23171
rect 18245 23137 18279 23171
rect 21465 23137 21499 23171
rect 24041 23137 24075 23171
rect 24961 23137 24995 23171
rect 5641 23069 5675 23103
rect 7849 23069 7883 23103
rect 10609 23069 10643 23103
rect 11437 23069 11471 23103
rect 12265 23069 12299 23103
rect 12633 23069 12667 23103
rect 12725 23069 12759 23103
rect 13277 23069 13311 23103
rect 13553 23069 13587 23103
rect 14473 23069 14507 23103
rect 14657 23069 14691 23103
rect 15833 23069 15867 23103
rect 17693 23069 17727 23103
rect 19349 23069 19383 23103
rect 21005 23069 21039 23103
rect 21189 23069 21223 23103
rect 21732 23069 21766 23103
rect 24685 23069 24719 23103
rect 5886 23001 5920 23035
rect 10342 23001 10376 23035
rect 11713 23001 11747 23035
rect 13001 23001 13035 23035
rect 14933 23001 14967 23035
rect 17969 23001 18003 23035
rect 19594 23001 19628 23035
rect 7021 22933 7055 22967
rect 8401 22933 8435 22967
rect 9229 22933 9263 22967
rect 11621 22933 11655 22967
rect 11805 22933 11839 22967
rect 13369 22933 13403 22967
rect 17785 22933 17819 22967
rect 18889 22933 18923 22967
rect 4629 22729 4663 22763
rect 8677 22729 8711 22763
rect 12633 22729 12667 22763
rect 14289 22729 14323 22763
rect 18521 22729 18555 22763
rect 19809 22729 19843 22763
rect 23765 22729 23799 22763
rect 24133 22729 24167 22763
rect 13746 22661 13780 22695
rect 18889 22661 18923 22695
rect 22652 22661 22686 22695
rect 4445 22593 4479 22627
rect 8401 22593 8435 22627
rect 8493 22593 8527 22627
rect 9413 22593 9447 22627
rect 9680 22593 9714 22627
rect 14841 22593 14875 22627
rect 18429 22593 18463 22627
rect 18521 22593 18555 22627
rect 19441 22593 19475 22627
rect 19993 22593 20027 22627
rect 20085 22593 20119 22627
rect 22385 22593 22419 22627
rect 24041 22593 24075 22627
rect 24225 22593 24259 22627
rect 4261 22525 4295 22559
rect 4997 22525 5031 22559
rect 12173 22525 12207 22559
rect 14013 22525 14047 22559
rect 18245 22525 18279 22559
rect 10793 22457 10827 22491
rect 9045 22389 9079 22423
rect 11161 22389 11195 22423
rect 11621 22389 11655 22423
rect 10701 22185 10735 22219
rect 12449 22185 12483 22219
rect 14841 22185 14875 22219
rect 18705 22185 18739 22219
rect 9781 22049 9815 22083
rect 10425 22049 10459 22083
rect 11069 22049 11103 22083
rect 23213 22049 23247 22083
rect 1501 21981 1535 22015
rect 1961 21981 1995 22015
rect 10885 21981 10919 22015
rect 11621 21981 11655 22015
rect 13829 21981 13863 22015
rect 14197 21981 14231 22015
rect 23121 21981 23155 22015
rect 23305 21981 23339 22015
rect 13562 21913 13596 21947
rect 17233 21913 17267 21947
rect 1685 21845 1719 21879
rect 12173 21845 12207 21879
rect 16865 21845 16899 21879
rect 12081 21641 12115 21675
rect 11621 21573 11655 21607
rect 10885 21505 10919 21539
rect 11069 21505 11103 21539
rect 11805 21505 11839 21539
rect 11897 21505 11931 21539
rect 12725 21505 12759 21539
rect 10425 21369 10459 21403
rect 10701 21301 10735 21335
rect 11897 21301 11931 21335
rect 12633 21301 12667 21335
rect 13093 21301 13127 21335
rect 11897 21097 11931 21131
rect 13553 21097 13587 21131
rect 10517 20961 10551 20995
rect 12173 20961 12207 20995
rect 10784 20893 10818 20927
rect 14933 20893 14967 20927
rect 15117 20893 15151 20927
rect 15577 20893 15611 20927
rect 12440 20825 12474 20859
rect 16221 20825 16255 20859
rect 15025 20757 15059 20791
rect 12449 20553 12483 20587
rect 14832 20485 14866 20519
rect 19809 20485 19843 20519
rect 20009 20485 20043 20519
rect 21925 20485 21959 20519
rect 22125 20485 22159 20519
rect 6469 20417 6503 20451
rect 6725 20417 6759 20451
rect 12173 20417 12207 20451
rect 12265 20417 12299 20451
rect 12725 20417 12759 20451
rect 21281 20417 21315 20451
rect 22569 20417 22603 20451
rect 22753 20417 22787 20451
rect 14565 20349 14599 20383
rect 21097 20349 21131 20383
rect 22293 20281 22327 20315
rect 7849 20213 7883 20247
rect 15945 20213 15979 20247
rect 19993 20213 20027 20247
rect 20177 20213 20211 20247
rect 21465 20213 21499 20247
rect 22109 20213 22143 20247
rect 22569 20213 22603 20247
rect 5641 20009 5675 20043
rect 6377 20009 6411 20043
rect 22477 20009 22511 20043
rect 23581 20009 23615 20043
rect 16221 19941 16255 19975
rect 17785 19941 17819 19975
rect 8125 19873 8159 19907
rect 14565 19873 14599 19907
rect 18245 19873 18279 19907
rect 22937 19873 22971 19907
rect 6101 19805 6135 19839
rect 6193 19805 6227 19839
rect 7297 19805 7331 19839
rect 16405 19805 16439 19839
rect 16497 19805 16531 19839
rect 17601 19805 17635 19839
rect 17877 19805 17911 19839
rect 18153 19805 18187 19839
rect 18331 19805 18365 19839
rect 18797 19805 18831 19839
rect 18889 19805 18923 19839
rect 19533 19805 19567 19839
rect 20821 19805 20855 19839
rect 21833 19805 21867 19839
rect 22753 19805 22787 19839
rect 6653 19737 6687 19771
rect 14832 19737 14866 19771
rect 16221 19737 16255 19771
rect 20177 19737 20211 19771
rect 7573 19669 7607 19703
rect 15945 19669 15979 19703
rect 17417 19669 17451 19703
rect 18613 19669 18647 19703
rect 21373 19669 21407 19703
rect 7849 19465 7883 19499
rect 13461 19465 13495 19499
rect 15025 19465 15059 19499
rect 19533 19465 19567 19499
rect 23305 19465 23339 19499
rect 24317 19465 24351 19499
rect 8984 19397 9018 19431
rect 10793 19397 10827 19431
rect 15761 19397 15795 19431
rect 5641 19329 5675 19363
rect 9229 19329 9263 19363
rect 10609 19329 10643 19363
rect 13553 19329 13587 19363
rect 15209 19329 15243 19363
rect 16037 19329 16071 19363
rect 16773 19329 16807 19363
rect 18420 19329 18454 19363
rect 19809 19329 19843 19363
rect 20729 19329 20763 19363
rect 21281 19329 21315 19363
rect 21925 19329 21959 19363
rect 22109 19329 22143 19363
rect 5825 19261 5859 19295
rect 6469 19261 6503 19295
rect 7113 19261 7147 19295
rect 10057 19261 10091 19295
rect 10425 19261 10459 19295
rect 15485 19261 15519 19295
rect 17325 19261 17359 19295
rect 18153 19261 18187 19295
rect 20361 19261 20395 19295
rect 22385 19261 22419 19295
rect 23857 19261 23891 19295
rect 15393 19193 15427 19227
rect 15945 19193 15979 19227
rect 5457 19125 5491 19159
rect 9505 19125 9539 19159
rect 15853 19125 15887 19159
rect 21925 19125 21959 19159
rect 23029 19125 23063 19159
rect 10517 18921 10551 18955
rect 18981 18921 19015 18955
rect 19441 18921 19475 18955
rect 19809 18921 19843 18955
rect 21741 18921 21775 18955
rect 23673 18853 23707 18887
rect 7481 18785 7515 18819
rect 10793 18785 10827 18819
rect 10885 18785 10919 18819
rect 11253 18785 11287 18819
rect 15117 18785 15151 18819
rect 19349 18785 19383 18819
rect 23397 18785 23431 18819
rect 24501 18785 24535 18819
rect 4077 18717 4111 18751
rect 4261 18717 4295 18751
rect 5273 18717 5307 18751
rect 7205 18717 7239 18751
rect 9045 18717 9079 18751
rect 9229 18717 9263 18751
rect 9413 18717 9447 18751
rect 9873 18717 9907 18751
rect 11161 18717 11195 18751
rect 15945 18717 15979 18751
rect 17601 18717 17635 18751
rect 19625 18717 19659 18751
rect 20361 18717 20395 18751
rect 23130 18717 23164 18751
rect 23673 18717 23707 18751
rect 23949 18717 23983 18751
rect 5540 18649 5574 18683
rect 6929 18649 6963 18683
rect 7297 18649 7331 18683
rect 7757 18649 7791 18683
rect 9321 18649 9355 18683
rect 11437 18649 11471 18683
rect 15669 18649 15703 18683
rect 16190 18649 16224 18683
rect 17846 18649 17880 18683
rect 20628 18649 20662 18683
rect 25145 18649 25179 18683
rect 4445 18581 4479 18615
rect 6653 18581 6687 18615
rect 7113 18581 7147 18615
rect 9597 18581 9631 18615
rect 10977 18581 11011 18615
rect 17325 18581 17359 18615
rect 22017 18581 22051 18615
rect 23857 18581 23891 18615
rect 3801 18377 3835 18411
rect 6101 18377 6135 18411
rect 7849 18377 7883 18411
rect 9413 18377 9447 18411
rect 15662 18377 15696 18411
rect 20821 18377 20855 18411
rect 22385 18377 22419 18411
rect 16205 18309 16239 18343
rect 16405 18309 16439 18343
rect 16773 18309 16807 18343
rect 4721 18241 4755 18275
rect 4988 18241 5022 18275
rect 6653 18241 6687 18275
rect 6745 18241 6779 18275
rect 6929 18241 6963 18275
rect 8125 18241 8159 18275
rect 11069 18241 11103 18275
rect 15485 18241 15519 18275
rect 15577 18241 15611 18275
rect 15761 18241 15795 18275
rect 17325 18241 17359 18275
rect 18613 18241 18647 18275
rect 21005 18241 21039 18275
rect 21189 18241 21223 18275
rect 21925 18241 21959 18275
rect 22017 18241 22051 18275
rect 22201 18241 22235 18275
rect 23785 18241 23819 18275
rect 24041 18241 24075 18275
rect 4445 18173 4479 18207
rect 7297 18173 7331 18207
rect 10701 18173 10735 18207
rect 12173 18173 12207 18207
rect 21281 18173 21315 18207
rect 6469 18105 6503 18139
rect 1501 18037 1535 18071
rect 6929 18037 6963 18071
rect 10149 18037 10183 18071
rect 11621 18037 11655 18071
rect 16037 18037 16071 18071
rect 16221 18037 16255 18071
rect 22661 18037 22695 18071
rect 6009 17833 6043 17867
rect 8217 17833 8251 17867
rect 11713 17833 11747 17867
rect 16773 17833 16807 17867
rect 21005 17833 21039 17867
rect 24501 17833 24535 17867
rect 24869 17833 24903 17867
rect 11345 17765 11379 17799
rect 19533 17765 19567 17799
rect 2973 17697 3007 17731
rect 9965 17697 9999 17731
rect 17325 17697 17359 17731
rect 19349 17697 19383 17731
rect 19809 17697 19843 17731
rect 23305 17697 23339 17731
rect 3157 17629 3191 17663
rect 4629 17629 4663 17663
rect 4896 17629 4930 17663
rect 6837 17629 6871 17663
rect 9321 17629 9355 17663
rect 9505 17629 9539 17663
rect 9689 17629 9723 17663
rect 11897 17629 11931 17663
rect 12173 17629 12207 17663
rect 15025 17629 15059 17663
rect 15117 17629 15151 17663
rect 15301 17629 15335 17663
rect 15393 17629 15427 17663
rect 15945 17629 15979 17663
rect 16313 17629 16347 17663
rect 17877 17629 17911 17663
rect 17970 17629 18004 17663
rect 18342 17629 18376 17663
rect 20177 17629 20211 17663
rect 20545 17629 20579 17663
rect 21005 17629 21039 17663
rect 21189 17629 21223 17663
rect 21557 17629 21591 17663
rect 21741 17629 21775 17663
rect 21833 17629 21867 17663
rect 21925 17629 21959 17663
rect 22109 17629 22143 17663
rect 24685 17629 24719 17663
rect 24961 17629 24995 17663
rect 7082 17561 7116 17595
rect 10210 17561 10244 17595
rect 15577 17561 15611 17595
rect 16129 17561 16163 17595
rect 16221 17561 16255 17595
rect 18153 17561 18187 17595
rect 18245 17561 18279 17595
rect 20361 17561 20395 17595
rect 20453 17561 20487 17595
rect 3341 17493 3375 17527
rect 16497 17493 16531 17527
rect 18521 17493 18555 17527
rect 20729 17493 20763 17527
rect 22293 17493 22327 17527
rect 23949 17493 23983 17527
rect 1685 17289 1719 17323
rect 5457 17289 5491 17323
rect 6101 17289 6135 17323
rect 7389 17289 7423 17323
rect 9505 17289 9539 17323
rect 11161 17289 11195 17323
rect 15853 17289 15887 17323
rect 17601 17289 17635 17323
rect 18061 17289 18095 17323
rect 20453 17289 20487 17323
rect 10048 17221 10082 17255
rect 15485 17221 15519 17255
rect 18429 17221 18463 17255
rect 1501 17153 1535 17187
rect 1961 17153 1995 17187
rect 3341 17153 3375 17187
rect 3597 17153 3631 17187
rect 5273 17153 5307 17187
rect 5825 17153 5859 17187
rect 5917 17153 5951 17187
rect 6745 17153 6779 17187
rect 8381 17153 8415 17187
rect 9781 17153 9815 17187
rect 12265 17153 12299 17187
rect 12449 17153 12483 17187
rect 15669 17153 15703 17187
rect 17049 17153 17083 17187
rect 17325 17153 17359 17187
rect 17417 17153 17451 17187
rect 20667 17153 20701 17187
rect 20821 17153 20855 17187
rect 22385 17153 22419 17187
rect 22569 17153 22603 17187
rect 23029 17153 23063 17187
rect 23121 17153 23155 17187
rect 23397 17153 23431 17187
rect 27261 17153 27295 17187
rect 5089 17085 5123 17119
rect 8125 17085 8159 17119
rect 17141 17085 17175 17119
rect 20177 17085 20211 17119
rect 22201 17085 22235 17119
rect 24317 17085 24351 17119
rect 28273 17085 28307 17119
rect 4721 16949 4755 16983
rect 12357 16949 12391 16983
rect 22845 16949 22879 16983
rect 23305 16949 23339 16983
rect 24961 16949 24995 16983
rect 7481 16745 7515 16779
rect 8125 16745 8159 16779
rect 23949 16745 23983 16779
rect 27537 16745 27571 16779
rect 6745 16609 6779 16643
rect 7757 16609 7791 16643
rect 8401 16609 8435 16643
rect 11805 16609 11839 16643
rect 12541 16609 12575 16643
rect 23857 16609 23891 16643
rect 24685 16609 24719 16643
rect 6101 16541 6135 16575
rect 7205 16541 7239 16575
rect 7297 16541 7331 16575
rect 7481 16541 7515 16575
rect 7941 16541 7975 16575
rect 12173 16541 12207 16575
rect 12449 16541 12483 16575
rect 12725 16541 12759 16575
rect 13277 16541 13311 16575
rect 23489 16541 23523 16575
rect 23765 16541 23799 16575
rect 24952 16541 24986 16575
rect 27721 16541 27755 16575
rect 27997 16541 28031 16575
rect 13093 16473 13127 16507
rect 7021 16405 7055 16439
rect 13461 16405 13495 16439
rect 23581 16405 23615 16439
rect 26065 16405 26099 16439
rect 14013 16201 14047 16235
rect 11805 16065 11839 16099
rect 12449 16065 12483 16099
rect 13185 16065 13219 16099
rect 13277 16065 13311 16099
rect 13921 16065 13955 16099
rect 14197 16065 14231 16099
rect 14657 16065 14691 16099
rect 27077 16065 27111 16099
rect 11897 15997 11931 16031
rect 28273 15997 28307 16031
rect 12173 15929 12207 15963
rect 12725 15929 12759 15963
rect 14381 15929 14415 15963
rect 14749 15861 14783 15895
rect 24041 15861 24075 15895
rect 12725 15657 12759 15691
rect 13645 15657 13679 15691
rect 14841 15657 14875 15691
rect 12081 15589 12115 15623
rect 13829 15589 13863 15623
rect 15209 15521 15243 15555
rect 10701 15453 10735 15487
rect 12357 15453 12391 15487
rect 12725 15453 12759 15487
rect 12909 15453 12943 15487
rect 14197 15453 14231 15487
rect 14657 15453 14691 15487
rect 15393 15453 15427 15487
rect 15761 15453 15795 15487
rect 10968 15385 11002 15419
rect 13461 15385 13495 15419
rect 15669 15385 15703 15419
rect 12541 15317 12575 15351
rect 13661 15317 13695 15351
rect 11621 15113 11655 15147
rect 14289 15113 14323 15147
rect 9321 14977 9355 15011
rect 11805 14977 11839 15011
rect 11897 14977 11931 15011
rect 15117 14977 15151 15011
rect 23765 14977 23799 15011
rect 13645 14909 13679 14943
rect 14381 14909 14415 14943
rect 14473 14909 14507 14943
rect 14933 14909 14967 14943
rect 24685 14909 24719 14943
rect 13921 14841 13955 14875
rect 13001 14773 13035 14807
rect 15301 14773 15335 14807
rect 23673 14773 23707 14807
rect 24041 14773 24075 14807
rect 8493 14569 8527 14603
rect 9781 14569 9815 14603
rect 11345 14569 11379 14603
rect 11989 14569 12023 14603
rect 13553 14569 13587 14603
rect 15117 14569 15151 14603
rect 25145 14569 25179 14603
rect 25421 14569 25455 14603
rect 8677 14501 8711 14535
rect 24133 14501 24167 14535
rect 12633 14433 12667 14467
rect 13369 14433 13403 14467
rect 15485 14433 15519 14467
rect 20729 14433 20763 14467
rect 22753 14433 22787 14467
rect 24501 14433 24535 14467
rect 7757 14365 7791 14399
rect 7941 14365 7975 14399
rect 8401 14365 8435 14399
rect 8493 14365 8527 14399
rect 11069 14365 11103 14399
rect 13277 14365 13311 14399
rect 14473 14365 14507 14399
rect 15393 14365 15427 14399
rect 15577 14365 15611 14399
rect 21005 14365 21039 14399
rect 25421 14365 25455 14399
rect 25605 14365 25639 14399
rect 28457 14365 28491 14399
rect 8217 14297 8251 14331
rect 20462 14297 20496 14331
rect 23020 14297 23054 14331
rect 7573 14229 7607 14263
rect 19349 14229 19383 14263
rect 21649 14229 21683 14263
rect 8769 14025 8803 14059
rect 14381 14025 14415 14059
rect 14749 14025 14783 14059
rect 20269 14025 20303 14059
rect 23213 14025 23247 14059
rect 9873 13957 9907 13991
rect 9965 13957 9999 13991
rect 10517 13957 10551 13991
rect 20637 13957 20671 13991
rect 9781 13889 9815 13923
rect 10149 13889 10183 13923
rect 13001 13889 13035 13923
rect 13268 13889 13302 13923
rect 14841 13889 14875 13923
rect 18981 13889 19015 13923
rect 19165 13889 19199 13923
rect 20545 13889 20579 13923
rect 20821 13889 20855 13923
rect 21097 13889 21131 13923
rect 24501 13889 24535 13923
rect 7481 13821 7515 13855
rect 8125 13821 8159 13855
rect 11161 13821 11195 13855
rect 18889 13821 18923 13855
rect 19349 13821 19383 13855
rect 19625 13821 19659 13855
rect 23765 13821 23799 13855
rect 24409 13821 24443 13855
rect 20821 13753 20855 13787
rect 6929 13685 6963 13719
rect 9597 13685 9631 13719
rect 24225 13685 24259 13719
rect 8125 13481 8159 13515
rect 10333 13481 10367 13515
rect 11989 13481 12023 13515
rect 13553 13481 13587 13515
rect 23581 13413 23615 13447
rect 10149 13345 10183 13379
rect 10609 13345 10643 13379
rect 16589 13345 16623 13379
rect 17509 13345 17543 13379
rect 20729 13345 20763 13379
rect 23121 13345 23155 13379
rect 6745 13277 6779 13311
rect 9137 13277 9171 13311
rect 9229 13277 9263 13311
rect 9689 13277 9723 13311
rect 10057 13277 10091 13311
rect 13553 13277 13587 13311
rect 13737 13277 13771 13311
rect 16681 13277 16715 13311
rect 17325 13277 17359 13311
rect 17417 13277 17451 13311
rect 17601 13277 17635 13311
rect 19901 13277 19935 13311
rect 20085 13277 20119 13311
rect 20269 13277 20303 13311
rect 20636 13277 20670 13311
rect 20821 13277 20855 13311
rect 20913 13277 20947 13311
rect 23213 13277 23247 13311
rect 7012 13209 7046 13243
rect 9413 13209 9447 13243
rect 9781 13209 9815 13243
rect 10876 13209 10910 13243
rect 19993 13209 20027 13243
rect 9965 13141 9999 13175
rect 14289 13141 14323 13175
rect 16313 13141 16347 13175
rect 17141 13141 17175 13175
rect 19717 13141 19751 13175
rect 21097 13141 21131 13175
rect 23857 13141 23891 13175
rect 7021 12937 7055 12971
rect 8677 12937 8711 12971
rect 9597 12937 9631 12971
rect 10885 12937 10919 12971
rect 13001 12937 13035 12971
rect 16405 12937 16439 12971
rect 17233 12937 17267 12971
rect 19809 12937 19843 12971
rect 22385 12937 22419 12971
rect 24133 12937 24167 12971
rect 24961 12937 24995 12971
rect 7564 12869 7598 12903
rect 12265 12869 12299 12903
rect 17877 12869 17911 12903
rect 23765 12869 23799 12903
rect 24225 12869 24259 12903
rect 5917 12801 5951 12835
rect 6745 12801 6779 12835
rect 6837 12801 6871 12835
rect 7297 12801 7331 12835
rect 8953 12801 8987 12835
rect 10241 12801 10275 12835
rect 12541 12801 12575 12835
rect 12817 12801 12851 12835
rect 16037 12801 16071 12835
rect 17141 12801 17175 12835
rect 17785 12801 17819 12835
rect 18061 12801 18095 12835
rect 18521 12801 18555 12835
rect 19441 12801 19475 12835
rect 20453 12801 20487 12835
rect 21281 12801 21315 12835
rect 22017 12801 22051 12835
rect 22201 12801 22235 12835
rect 23121 12801 23155 12835
rect 23857 12801 23891 12835
rect 23949 12801 23983 12835
rect 24501 12801 24535 12835
rect 24593 12801 24627 12835
rect 24777 12801 24811 12835
rect 6101 12733 6135 12767
rect 11621 12733 11655 12767
rect 12633 12733 12667 12767
rect 16129 12733 16163 12767
rect 17417 12733 17451 12767
rect 19349 12733 19383 12767
rect 20085 12733 20119 12767
rect 20361 12733 20395 12767
rect 21189 12733 21223 12767
rect 21925 12733 21959 12767
rect 23029 12733 23063 12767
rect 18613 12665 18647 12699
rect 20913 12665 20947 12699
rect 23489 12665 23523 12699
rect 5733 12597 5767 12631
rect 12541 12597 12575 12631
rect 16773 12597 16807 12631
rect 18245 12597 18279 12631
rect 11345 12393 11379 12427
rect 11621 12393 11655 12427
rect 18337 12393 18371 12427
rect 8677 12325 8711 12359
rect 18613 12325 18647 12359
rect 23857 12325 23891 12359
rect 9137 12257 9171 12291
rect 15761 12257 15795 12291
rect 16865 12257 16899 12291
rect 18981 12257 19015 12291
rect 19717 12257 19751 12291
rect 20821 12257 20855 12291
rect 23305 12257 23339 12291
rect 23397 12257 23431 12291
rect 24501 12257 24535 12291
rect 5641 12189 5675 12223
rect 7297 12189 7331 12223
rect 9965 12189 9999 12223
rect 13001 12189 13035 12223
rect 15669 12189 15703 12223
rect 17785 12189 17819 12223
rect 18797 12189 18831 12223
rect 19625 12189 19659 12223
rect 21833 12189 21867 12223
rect 22753 12189 22787 12223
rect 5886 12121 5920 12155
rect 7564 12121 7598 12155
rect 10232 12121 10266 12155
rect 12734 12121 12768 12155
rect 20729 12121 20763 12155
rect 23489 12121 23523 12155
rect 7021 12053 7055 12087
rect 9689 12053 9723 12087
rect 16037 12053 16071 12087
rect 16313 12053 16347 12087
rect 19993 12053 20027 12087
rect 20269 12053 20303 12087
rect 20637 12053 20671 12087
rect 21281 12053 21315 12087
rect 22201 12053 22235 12087
rect 25145 12053 25179 12087
rect 6469 11849 6503 11883
rect 8585 11849 8619 11883
rect 16773 11849 16807 11883
rect 17601 11849 17635 11883
rect 21005 11849 21039 11883
rect 22477 11849 22511 11883
rect 22753 11849 22787 11883
rect 24869 11849 24903 11883
rect 21373 11781 21407 11815
rect 22017 11781 22051 11815
rect 23888 11781 23922 11815
rect 25237 11781 25271 11815
rect 5549 11713 5583 11747
rect 5641 11713 5675 11747
rect 8309 11713 8343 11747
rect 9709 11713 9743 11747
rect 9965 11713 9999 11747
rect 11253 11713 11287 11747
rect 14381 11713 14415 11747
rect 14565 11713 14599 11747
rect 15669 11713 15703 11747
rect 15853 11713 15887 11747
rect 17141 11713 17175 11747
rect 17785 11713 17819 11747
rect 19892 11713 19926 11747
rect 21465 11713 21499 11747
rect 24133 11713 24167 11747
rect 24685 11713 24719 11747
rect 25145 11713 25179 11747
rect 25329 11713 25363 11747
rect 25605 11713 25639 11747
rect 7113 11645 7147 11679
rect 14657 11645 14691 11679
rect 16129 11645 16163 11679
rect 17049 11645 17083 11679
rect 18061 11645 18095 11679
rect 19625 11645 19659 11679
rect 24501 11645 24535 11679
rect 22385 11577 22419 11611
rect 5825 11509 5859 11543
rect 7665 11509 7699 11543
rect 10609 11509 10643 11543
rect 14197 11509 14231 11543
rect 15853 11509 15887 11543
rect 17969 11509 18003 11543
rect 6837 11305 6871 11339
rect 7941 11305 7975 11339
rect 9597 11305 9631 11339
rect 10609 11305 10643 11339
rect 14933 11305 14967 11339
rect 16773 11305 16807 11339
rect 18153 11305 18187 11339
rect 19901 11305 19935 11339
rect 22109 11305 22143 11339
rect 22477 11305 22511 11339
rect 23857 11305 23891 11339
rect 9045 11237 9079 11271
rect 13829 11237 13863 11271
rect 23489 11237 23523 11271
rect 24501 11237 24535 11271
rect 5457 11169 5491 11203
rect 8309 11169 8343 11203
rect 10241 11169 10275 11203
rect 12449 11169 12483 11203
rect 14289 11169 14323 11203
rect 17509 11169 17543 11203
rect 17601 11169 17635 11203
rect 20729 11169 20763 11203
rect 5724 11101 5758 11135
rect 8125 11101 8159 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 10425 11101 10459 11135
rect 15393 11101 15427 11135
rect 18245 11101 18279 11135
rect 19717 11101 19751 11135
rect 19901 11101 19935 11135
rect 20177 11101 20211 11135
rect 21741 11101 21775 11135
rect 21925 11101 21959 11135
rect 22569 11101 22603 11135
rect 9229 11033 9263 11067
rect 12716 11033 12750 11067
rect 15660 11033 15694 11067
rect 17417 11033 17451 11067
rect 23213 11033 23247 11067
rect 17049 10965 17083 10999
rect 9505 10761 9539 10795
rect 13461 10761 13495 10795
rect 14565 10761 14599 10795
rect 18521 10761 18555 10795
rect 19993 10761 20027 10795
rect 14381 10693 14415 10727
rect 15025 10693 15059 10727
rect 9689 10625 9723 10659
rect 9873 10625 9907 10659
rect 14105 10625 14139 10659
rect 14657 10625 14691 10659
rect 17325 10625 17359 10659
rect 17877 10625 17911 10659
rect 14381 10489 14415 10523
rect 16773 10421 16807 10455
rect 17601 10217 17635 10251
rect 16221 10081 16255 10115
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 15853 9945 15887 9979
rect 16466 9945 16500 9979
rect 16037 9673 16071 9707
rect 28273 8585 28307 8619
rect 27905 8449 27939 8483
rect 28457 8449 28491 8483
rect 28365 8041 28399 8075
rect 5917 2601 5951 2635
rect 6101 2397 6135 2431
rect 6469 2397 6503 2431
rect 22017 2397 22051 2431
<< metal1 >>
rect 1104 47354 28888 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 28888 47354
rect 1104 47280 28888 47302
rect 24578 47200 24584 47252
rect 24636 47200 24642 47252
rect 4706 47132 4712 47184
rect 4764 47172 4770 47184
rect 5261 47175 5319 47181
rect 5261 47172 5273 47175
rect 4764 47144 5273 47172
rect 4764 47132 4770 47144
rect 5261 47141 5273 47144
rect 5307 47141 5319 47175
rect 5261 47135 5319 47141
rect 22002 47064 22008 47116
rect 22060 47104 22066 47116
rect 22465 47107 22523 47113
rect 22465 47104 22477 47107
rect 22060 47076 22477 47104
rect 22060 47064 22066 47076
rect 22465 47073 22477 47076
rect 22511 47073 22523 47107
rect 22465 47067 22523 47073
rect 5442 46996 5448 47048
rect 5500 47036 5506 47048
rect 5721 47039 5779 47045
rect 5721 47036 5733 47039
rect 5500 47008 5733 47036
rect 5500 46996 5506 47008
rect 5721 47005 5733 47008
rect 5767 47005 5779 47039
rect 5721 46999 5779 47005
rect 22094 46996 22100 47048
rect 22152 46996 22158 47048
rect 1104 46810 28888 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 28888 46810
rect 1104 46736 28888 46758
rect 1104 46266 28888 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 28888 46266
rect 1104 46192 28888 46214
rect 1104 45722 28888 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 28888 45722
rect 1104 45648 28888 45670
rect 10042 45500 10048 45552
rect 10100 45540 10106 45552
rect 20622 45540 20628 45552
rect 10100 45512 12434 45540
rect 10100 45500 10106 45512
rect 10689 45475 10747 45481
rect 10689 45441 10701 45475
rect 10735 45441 10747 45475
rect 10689 45435 10747 45441
rect 10704 45404 10732 45435
rect 10870 45432 10876 45484
rect 10928 45432 10934 45484
rect 10980 45481 11008 45512
rect 10965 45475 11023 45481
rect 10965 45441 10977 45475
rect 11011 45441 11023 45475
rect 10965 45435 11023 45441
rect 11790 45432 11796 45484
rect 11848 45432 11854 45484
rect 11882 45432 11888 45484
rect 11940 45472 11946 45484
rect 11977 45475 12035 45481
rect 11977 45472 11989 45475
rect 11940 45444 11989 45472
rect 11940 45432 11946 45444
rect 11977 45441 11989 45444
rect 12023 45441 12035 45475
rect 11977 45435 12035 45441
rect 11698 45404 11704 45416
rect 10704 45376 11704 45404
rect 11698 45364 11704 45376
rect 11756 45364 11762 45416
rect 9950 45296 9956 45348
rect 10008 45336 10014 45348
rect 10870 45336 10876 45348
rect 10008 45308 10876 45336
rect 10008 45296 10014 45308
rect 10870 45296 10876 45308
rect 10928 45296 10934 45348
rect 12406 45336 12434 45512
rect 13924 45512 16068 45540
rect 13924 45484 13952 45512
rect 16040 45484 16068 45512
rect 17144 45512 20628 45540
rect 13817 45475 13875 45481
rect 13817 45441 13829 45475
rect 13863 45441 13875 45475
rect 13817 45435 13875 45441
rect 13832 45404 13860 45435
rect 13906 45432 13912 45484
rect 13964 45432 13970 45484
rect 14461 45475 14519 45481
rect 14461 45441 14473 45475
rect 14507 45441 14519 45475
rect 14461 45435 14519 45441
rect 14645 45475 14703 45481
rect 14645 45441 14657 45475
rect 14691 45472 14703 45475
rect 14734 45472 14740 45484
rect 14691 45444 14740 45472
rect 14691 45441 14703 45444
rect 14645 45435 14703 45441
rect 14366 45404 14372 45416
rect 13832 45376 14372 45404
rect 14366 45364 14372 45376
rect 14424 45364 14430 45416
rect 14476 45404 14504 45435
rect 14734 45432 14740 45444
rect 14792 45432 14798 45484
rect 16022 45432 16028 45484
rect 16080 45432 16086 45484
rect 17144 45481 17172 45512
rect 20622 45500 20628 45512
rect 20680 45500 20686 45552
rect 17129 45475 17187 45481
rect 17129 45441 17141 45475
rect 17175 45441 17187 45475
rect 17129 45435 17187 45441
rect 17313 45475 17371 45481
rect 17313 45441 17325 45475
rect 17359 45472 17371 45475
rect 19518 45472 19524 45484
rect 17359 45444 19524 45472
rect 17359 45441 17371 45444
rect 17313 45435 17371 45441
rect 19518 45432 19524 45444
rect 19576 45432 19582 45484
rect 19696 45475 19754 45481
rect 19696 45441 19708 45475
rect 19742 45472 19754 45475
rect 19978 45472 19984 45484
rect 19742 45444 19984 45472
rect 19742 45441 19754 45444
rect 19696 45435 19754 45441
rect 19978 45432 19984 45444
rect 20036 45432 20042 45484
rect 14476 45376 14964 45404
rect 14090 45336 14096 45348
rect 12406 45308 14096 45336
rect 14090 45296 14096 45308
rect 14148 45296 14154 45348
rect 14936 45280 14964 45376
rect 15746 45364 15752 45416
rect 15804 45404 15810 45416
rect 17037 45407 17095 45413
rect 17037 45404 17049 45407
rect 15804 45376 17049 45404
rect 15804 45364 15810 45376
rect 17037 45373 17049 45376
rect 17083 45404 17095 45407
rect 17083 45376 17816 45404
rect 17083 45373 17095 45376
rect 17037 45367 17095 45373
rect 17788 45280 17816 45376
rect 18138 45364 18144 45416
rect 18196 45404 18202 45416
rect 18325 45407 18383 45413
rect 18325 45404 18337 45407
rect 18196 45376 18337 45404
rect 18196 45364 18202 45376
rect 18325 45373 18337 45376
rect 18371 45373 18383 45407
rect 18325 45367 18383 45373
rect 18414 45364 18420 45416
rect 18472 45404 18478 45416
rect 19429 45407 19487 45413
rect 19429 45404 19441 45407
rect 18472 45376 19441 45404
rect 18472 45364 18478 45376
rect 19429 45373 19441 45376
rect 19475 45373 19487 45407
rect 19429 45367 19487 45373
rect 20809 45339 20867 45345
rect 20809 45305 20821 45339
rect 20855 45336 20867 45339
rect 22094 45336 22100 45348
rect 20855 45308 22100 45336
rect 20855 45305 20867 45308
rect 20809 45299 20867 45305
rect 22094 45296 22100 45308
rect 22152 45296 22158 45348
rect 9398 45228 9404 45280
rect 9456 45268 9462 45280
rect 10505 45271 10563 45277
rect 10505 45268 10517 45271
rect 9456 45240 10517 45268
rect 9456 45228 9462 45240
rect 10505 45237 10517 45240
rect 10551 45237 10563 45271
rect 10505 45231 10563 45237
rect 11054 45228 11060 45280
rect 11112 45268 11118 45280
rect 11609 45271 11667 45277
rect 11609 45268 11621 45271
rect 11112 45240 11621 45268
rect 11112 45228 11118 45240
rect 11609 45237 11621 45240
rect 11655 45237 11667 45271
rect 11609 45231 11667 45237
rect 13633 45271 13691 45277
rect 13633 45237 13645 45271
rect 13679 45268 13691 45271
rect 13814 45268 13820 45280
rect 13679 45240 13820 45268
rect 13679 45237 13691 45240
rect 13633 45231 13691 45237
rect 13814 45228 13820 45240
rect 13872 45228 13878 45280
rect 14642 45228 14648 45280
rect 14700 45228 14706 45280
rect 14918 45228 14924 45280
rect 14976 45228 14982 45280
rect 15933 45271 15991 45277
rect 15933 45237 15945 45271
rect 15979 45268 15991 45271
rect 16482 45268 16488 45280
rect 15979 45240 16488 45268
rect 15979 45237 15991 45240
rect 15933 45231 15991 45237
rect 16482 45228 16488 45240
rect 16540 45228 16546 45280
rect 17494 45228 17500 45280
rect 17552 45228 17558 45280
rect 17770 45228 17776 45280
rect 17828 45228 17834 45280
rect 1104 45178 28888 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 28888 45178
rect 1104 45104 28888 45126
rect 10042 45024 10048 45076
rect 10100 45024 10106 45076
rect 11698 45064 11704 45076
rect 10152 45036 11704 45064
rect 7466 44820 7472 44872
rect 7524 44820 7530 44872
rect 8021 44863 8079 44869
rect 8021 44829 8033 44863
rect 8067 44829 8079 44863
rect 8021 44823 8079 44829
rect 8205 44863 8263 44869
rect 8205 44829 8217 44863
rect 8251 44860 8263 44863
rect 9490 44860 9496 44872
rect 8251 44832 9496 44860
rect 8251 44829 8263 44832
rect 8205 44823 8263 44829
rect 8036 44792 8064 44823
rect 9490 44820 9496 44832
rect 9548 44820 9554 44872
rect 9861 44795 9919 44801
rect 8036 44764 8616 44792
rect 6914 44684 6920 44736
rect 6972 44684 6978 44736
rect 7834 44684 7840 44736
rect 7892 44684 7898 44736
rect 8588 44733 8616 44764
rect 9861 44761 9873 44795
rect 9907 44792 9919 44795
rect 9950 44792 9956 44804
rect 9907 44764 9956 44792
rect 9907 44761 9919 44764
rect 9861 44755 9919 44761
rect 9950 44752 9956 44764
rect 10008 44752 10014 44804
rect 10066 44795 10124 44801
rect 10066 44761 10078 44795
rect 10112 44792 10124 44795
rect 10152 44792 10180 45036
rect 11698 45024 11704 45036
rect 11756 45024 11762 45076
rect 16022 45024 16028 45076
rect 16080 45064 16086 45076
rect 16485 45067 16543 45073
rect 16485 45064 16497 45067
rect 16080 45036 16497 45064
rect 16080 45024 16086 45036
rect 16485 45033 16497 45036
rect 16531 45033 16543 45067
rect 16485 45027 16543 45033
rect 19978 45024 19984 45076
rect 20036 45024 20042 45076
rect 10229 44999 10287 45005
rect 10229 44965 10241 44999
rect 10275 44965 10287 44999
rect 10229 44959 10287 44965
rect 11241 44999 11299 45005
rect 11241 44965 11253 44999
rect 11287 44996 11299 44999
rect 15565 44999 15623 45005
rect 11287 44968 13032 44996
rect 11287 44965 11299 44968
rect 11241 44959 11299 44965
rect 10244 44928 10272 44959
rect 10873 44931 10931 44937
rect 10244 44900 10732 44928
rect 10704 44869 10732 44900
rect 10873 44897 10885 44931
rect 10919 44928 10931 44931
rect 11146 44928 11152 44940
rect 10919 44900 11152 44928
rect 10919 44897 10931 44900
rect 10873 44891 10931 44897
rect 11146 44888 11152 44900
rect 11204 44888 11210 44940
rect 13004 44937 13032 44968
rect 15565 44965 15577 44999
rect 15611 44996 15623 44999
rect 15611 44968 15884 44996
rect 15611 44965 15623 44968
rect 15565 44959 15623 44965
rect 15856 44937 15884 44968
rect 12989 44931 13047 44937
rect 12989 44897 13001 44931
rect 13035 44897 13047 44931
rect 12989 44891 13047 44897
rect 15841 44931 15899 44937
rect 15841 44897 15853 44931
rect 15887 44897 15899 44931
rect 15841 44891 15899 44897
rect 10505 44863 10563 44869
rect 10505 44829 10517 44863
rect 10551 44829 10563 44863
rect 10505 44823 10563 44829
rect 10689 44863 10747 44869
rect 10689 44829 10701 44863
rect 10735 44829 10747 44863
rect 10689 44823 10747 44829
rect 10112 44764 10180 44792
rect 10112 44761 10124 44764
rect 10066 44755 10124 44761
rect 8573 44727 8631 44733
rect 8573 44693 8585 44727
rect 8619 44724 8631 44727
rect 9214 44724 9220 44736
rect 8619 44696 9220 44724
rect 8619 44693 8631 44696
rect 8573 44687 8631 44693
rect 9214 44684 9220 44696
rect 9272 44684 9278 44736
rect 10520 44724 10548 44823
rect 10778 44820 10784 44872
rect 10836 44820 10842 44872
rect 11057 44863 11115 44869
rect 11057 44829 11069 44863
rect 11103 44829 11115 44863
rect 11057 44823 11115 44829
rect 11072 44792 11100 44823
rect 11238 44820 11244 44872
rect 11296 44860 11302 44872
rect 11517 44863 11575 44869
rect 11517 44860 11529 44863
rect 11296 44832 11529 44860
rect 11296 44820 11302 44832
rect 11517 44829 11529 44832
rect 11563 44829 11575 44863
rect 11517 44823 11575 44829
rect 11882 44820 11888 44872
rect 11940 44860 11946 44872
rect 14185 44863 14243 44869
rect 11940 44832 14136 44860
rect 11940 44820 11946 44832
rect 12161 44795 12219 44801
rect 12161 44792 12173 44795
rect 11072 44764 12173 44792
rect 12161 44761 12173 44764
rect 12207 44792 12219 44795
rect 12526 44792 12532 44804
rect 12207 44764 12532 44792
rect 12207 44761 12219 44764
rect 12161 44755 12219 44761
rect 12526 44752 12532 44764
rect 12584 44752 12590 44804
rect 14108 44792 14136 44832
rect 14185 44829 14197 44863
rect 14231 44860 14243 44863
rect 15010 44860 15016 44872
rect 14231 44832 15016 44860
rect 14231 44829 14243 44832
rect 14185 44823 14243 44829
rect 15010 44820 15016 44832
rect 15068 44860 15074 44872
rect 17129 44863 17187 44869
rect 17129 44860 17141 44863
rect 15068 44832 15240 44860
rect 15068 44820 15074 44832
rect 14274 44792 14280 44804
rect 14108 44764 14280 44792
rect 14274 44752 14280 44764
rect 14332 44752 14338 44804
rect 14452 44795 14510 44801
rect 14452 44761 14464 44795
rect 14498 44792 14510 44795
rect 14642 44792 14648 44804
rect 14498 44764 14648 44792
rect 14498 44761 14510 44764
rect 14452 44755 14510 44761
rect 14642 44752 14648 44764
rect 14700 44752 14706 44804
rect 15212 44792 15240 44832
rect 16546 44832 17141 44860
rect 16546 44792 16574 44832
rect 17129 44829 17141 44832
rect 17175 44860 17187 44863
rect 18414 44860 18420 44872
rect 17175 44832 18420 44860
rect 17175 44829 17187 44832
rect 17129 44823 17187 44829
rect 18414 44820 18420 44832
rect 18472 44820 18478 44872
rect 19334 44820 19340 44872
rect 19392 44820 19398 44872
rect 15212 44764 16574 44792
rect 17396 44795 17454 44801
rect 17396 44761 17408 44795
rect 17442 44792 17454 44795
rect 17494 44792 17500 44804
rect 17442 44764 17500 44792
rect 17442 44761 17454 44764
rect 17396 44755 17454 44761
rect 17494 44752 17500 44764
rect 17552 44752 17558 44804
rect 12250 44724 12256 44736
rect 10520 44696 12256 44724
rect 12250 44684 12256 44696
rect 12308 44684 12314 44736
rect 12434 44684 12440 44736
rect 12492 44684 12498 44736
rect 18138 44684 18144 44736
rect 18196 44724 18202 44736
rect 18509 44727 18567 44733
rect 18509 44724 18521 44727
rect 18196 44696 18521 44724
rect 18196 44684 18202 44696
rect 18509 44693 18521 44696
rect 18555 44693 18567 44727
rect 18509 44687 18567 44693
rect 1104 44634 28888 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 28888 44634
rect 1104 44560 28888 44582
rect 9585 44523 9643 44529
rect 9585 44489 9597 44523
rect 9631 44520 9643 44523
rect 10778 44520 10784 44532
rect 9631 44492 10784 44520
rect 9631 44489 9643 44492
rect 9585 44483 9643 44489
rect 10778 44480 10784 44492
rect 10836 44480 10842 44532
rect 11238 44480 11244 44532
rect 11296 44480 11302 44532
rect 11790 44480 11796 44532
rect 11848 44520 11854 44532
rect 11848 44492 13952 44520
rect 11848 44480 11854 44492
rect 6917 44455 6975 44461
rect 6917 44421 6929 44455
rect 6963 44452 6975 44455
rect 7438 44455 7496 44461
rect 7438 44452 7450 44455
rect 6963 44424 7450 44452
rect 6963 44421 6975 44424
rect 6917 44415 6975 44421
rect 7438 44421 7450 44424
rect 7484 44421 7496 44455
rect 7438 44415 7496 44421
rect 10128 44455 10186 44461
rect 10128 44421 10140 44455
rect 10174 44452 10186 44455
rect 12434 44452 12440 44464
rect 10174 44424 12440 44452
rect 10174 44421 10186 44424
rect 10128 44415 10186 44421
rect 12434 44412 12440 44424
rect 12492 44412 12498 44464
rect 13814 44452 13820 44464
rect 12820 44424 13820 44452
rect 4706 44344 4712 44396
rect 4764 44344 4770 44396
rect 4893 44387 4951 44393
rect 4893 44353 4905 44387
rect 4939 44384 4951 44387
rect 5626 44384 5632 44396
rect 4939 44356 5632 44384
rect 4939 44353 4951 44356
rect 4893 44347 4951 44353
rect 5626 44344 5632 44356
rect 5684 44384 5690 44396
rect 6733 44387 6791 44393
rect 6733 44384 6745 44387
rect 5684 44356 6745 44384
rect 5684 44344 5690 44356
rect 6733 44353 6745 44356
rect 6779 44353 6791 44387
rect 6733 44347 6791 44353
rect 9398 44344 9404 44396
rect 9456 44344 9462 44396
rect 9585 44387 9643 44393
rect 9585 44353 9597 44387
rect 9631 44384 9643 44387
rect 11146 44384 11152 44396
rect 9631 44356 11152 44384
rect 9631 44353 9643 44356
rect 9585 44347 9643 44353
rect 11146 44344 11152 44356
rect 11204 44344 11210 44396
rect 12529 44387 12587 44393
rect 12529 44384 12541 44387
rect 11624 44356 12541 44384
rect 6549 44319 6607 44325
rect 6549 44285 6561 44319
rect 6595 44285 6607 44319
rect 6549 44279 6607 44285
rect 4525 44183 4583 44189
rect 4525 44149 4537 44183
rect 4571 44180 4583 44183
rect 4706 44180 4712 44192
rect 4571 44152 4712 44180
rect 4571 44149 4583 44152
rect 4525 44143 4583 44149
rect 4706 44140 4712 44152
rect 4764 44140 4770 44192
rect 6564 44180 6592 44279
rect 7190 44276 7196 44328
rect 7248 44276 7254 44328
rect 9858 44276 9864 44328
rect 9916 44276 9922 44328
rect 11624 44325 11652 44356
rect 12529 44353 12541 44356
rect 12575 44353 12587 44387
rect 12529 44347 12587 44353
rect 12621 44387 12679 44393
rect 12621 44353 12633 44387
rect 12667 44384 12679 44387
rect 12710 44384 12716 44396
rect 12667 44356 12716 44384
rect 12667 44353 12679 44356
rect 12621 44347 12679 44353
rect 11609 44319 11667 44325
rect 11609 44285 11621 44319
rect 11655 44285 11667 44319
rect 11609 44279 11667 44285
rect 11698 44276 11704 44328
rect 11756 44316 11762 44328
rect 11793 44319 11851 44325
rect 11793 44316 11805 44319
rect 11756 44288 11805 44316
rect 11756 44276 11762 44288
rect 11793 44285 11805 44288
rect 11839 44285 11851 44319
rect 11793 44279 11851 44285
rect 11882 44276 11888 44328
rect 11940 44276 11946 44328
rect 11977 44319 12035 44325
rect 11977 44285 11989 44319
rect 12023 44285 12035 44319
rect 11977 44279 12035 44285
rect 12069 44319 12127 44325
rect 12069 44285 12081 44319
rect 12115 44316 12127 44319
rect 12115 44288 12434 44316
rect 12115 44285 12127 44288
rect 12069 44279 12127 44285
rect 11514 44208 11520 44260
rect 11572 44248 11578 44260
rect 11900 44248 11928 44276
rect 11572 44220 11928 44248
rect 11572 44208 11578 44220
rect 6914 44180 6920 44192
rect 6564 44152 6920 44180
rect 6914 44140 6920 44152
rect 6972 44180 6978 44192
rect 7926 44180 7932 44192
rect 6972 44152 7932 44180
rect 6972 44140 6978 44152
rect 7926 44140 7932 44152
rect 7984 44140 7990 44192
rect 8570 44140 8576 44192
rect 8628 44140 8634 44192
rect 11790 44140 11796 44192
rect 11848 44180 11854 44192
rect 11992 44180 12020 44279
rect 11848 44152 12020 44180
rect 12406 44180 12434 44288
rect 12544 44248 12572 44347
rect 12710 44344 12716 44356
rect 12768 44344 12774 44396
rect 12820 44393 12848 44424
rect 13814 44412 13820 44424
rect 13872 44412 13878 44464
rect 12805 44387 12863 44393
rect 12805 44353 12817 44387
rect 12851 44353 12863 44387
rect 12805 44347 12863 44353
rect 13446 44344 13452 44396
rect 13504 44344 13510 44396
rect 13924 44384 13952 44492
rect 14090 44480 14096 44532
rect 14148 44480 14154 44532
rect 14645 44523 14703 44529
rect 14645 44489 14657 44523
rect 14691 44520 14703 44523
rect 14734 44520 14740 44532
rect 14691 44492 14740 44520
rect 14691 44489 14703 44492
rect 14645 44483 14703 44489
rect 14734 44480 14740 44492
rect 14792 44480 14798 44532
rect 17770 44480 17776 44532
rect 17828 44520 17834 44532
rect 20533 44523 20591 44529
rect 20533 44520 20545 44523
rect 17828 44492 20545 44520
rect 17828 44480 17834 44492
rect 20533 44489 20545 44492
rect 20579 44489 20591 44523
rect 20533 44483 20591 44489
rect 15013 44455 15071 44461
rect 15013 44421 15025 44455
rect 15059 44452 15071 44455
rect 16482 44452 16488 44464
rect 15059 44424 16488 44452
rect 15059 44421 15071 44424
rect 15013 44415 15071 44421
rect 16482 44412 16488 44424
rect 16540 44412 16546 44464
rect 18230 44452 18236 44464
rect 17788 44424 18236 44452
rect 14093 44387 14151 44393
rect 14093 44384 14105 44387
rect 13924 44356 14105 44384
rect 14093 44353 14105 44356
rect 14139 44353 14151 44387
rect 14093 44347 14151 44353
rect 14274 44344 14280 44396
rect 14332 44344 14338 44396
rect 15746 44344 15752 44396
rect 15804 44384 15810 44396
rect 17788 44393 17816 44424
rect 18230 44412 18236 44424
rect 18288 44452 18294 44464
rect 18414 44452 18420 44464
rect 18288 44424 18420 44452
rect 18288 44412 18294 44424
rect 18414 44412 18420 44424
rect 18472 44412 18478 44464
rect 18046 44393 18052 44396
rect 16025 44387 16083 44393
rect 16025 44384 16037 44387
rect 15804 44356 16037 44384
rect 15804 44344 15810 44356
rect 16025 44353 16037 44356
rect 16071 44353 16083 44387
rect 16025 44347 16083 44353
rect 16118 44387 16176 44393
rect 16118 44353 16130 44387
rect 16164 44384 16176 44387
rect 16761 44387 16819 44393
rect 16761 44384 16773 44387
rect 16164 44356 16773 44384
rect 16164 44353 16176 44356
rect 16118 44347 16176 44353
rect 16761 44353 16773 44356
rect 16807 44353 16819 44387
rect 16761 44347 16819 44353
rect 17773 44387 17831 44393
rect 17773 44353 17785 44387
rect 17819 44353 17831 44387
rect 17773 44347 17831 44353
rect 18040 44347 18052 44393
rect 13357 44319 13415 44325
rect 13357 44285 13369 44319
rect 13403 44285 13415 44319
rect 15105 44319 15163 44325
rect 15105 44316 15117 44319
rect 13357 44279 13415 44285
rect 13832 44288 15117 44316
rect 13372 44248 13400 44279
rect 13832 44257 13860 44288
rect 15105 44285 15117 44288
rect 15151 44285 15163 44319
rect 15105 44279 15163 44285
rect 15197 44319 15255 44325
rect 15197 44285 15209 44319
rect 15243 44285 15255 44319
rect 15197 44279 15255 44285
rect 12544 44220 13400 44248
rect 13817 44251 13875 44257
rect 13817 44217 13829 44251
rect 13863 44217 13875 44251
rect 13817 44211 13875 44217
rect 14734 44208 14740 44260
rect 14792 44248 14798 44260
rect 15212 44248 15240 44279
rect 15562 44276 15568 44328
rect 15620 44316 15626 44328
rect 16132 44316 16160 44347
rect 18046 44344 18052 44347
rect 18104 44344 18110 44396
rect 20349 44387 20407 44393
rect 20349 44353 20361 44387
rect 20395 44353 20407 44387
rect 20349 44347 20407 44353
rect 15620 44288 16160 44316
rect 15620 44276 15626 44288
rect 16850 44276 16856 44328
rect 16908 44316 16914 44328
rect 17313 44319 17371 44325
rect 17313 44316 17325 44319
rect 16908 44288 17325 44316
rect 16908 44276 16914 44288
rect 17313 44285 17325 44288
rect 17359 44285 17371 44319
rect 17313 44279 17371 44285
rect 19429 44319 19487 44325
rect 19429 44285 19441 44319
rect 19475 44285 19487 44319
rect 20364 44316 20392 44347
rect 20622 44344 20628 44396
rect 20680 44344 20686 44396
rect 20364 44288 21036 44316
rect 19429 44279 19487 44285
rect 14792 44220 15240 44248
rect 16393 44251 16451 44257
rect 14792 44208 14798 44220
rect 16393 44217 16405 44251
rect 16439 44248 16451 44251
rect 17678 44248 17684 44260
rect 16439 44220 17684 44248
rect 16439 44217 16451 44220
rect 16393 44211 16451 44217
rect 17678 44208 17684 44220
rect 17736 44208 17742 44260
rect 19153 44251 19211 44257
rect 19153 44217 19165 44251
rect 19199 44248 19211 44251
rect 19444 44248 19472 44279
rect 19199 44220 19472 44248
rect 19199 44217 19211 44220
rect 19153 44211 19211 44217
rect 19518 44208 19524 44260
rect 19576 44248 19582 44260
rect 20349 44251 20407 44257
rect 20349 44248 20361 44251
rect 19576 44220 20361 44248
rect 19576 44208 19582 44220
rect 20349 44217 20361 44220
rect 20395 44217 20407 44251
rect 20349 44211 20407 44217
rect 12894 44180 12900 44192
rect 12406 44152 12900 44180
rect 11848 44140 11854 44152
rect 12894 44140 12900 44152
rect 12952 44140 12958 44192
rect 12989 44183 13047 44189
rect 12989 44149 13001 44183
rect 13035 44180 13047 44183
rect 13998 44180 14004 44192
rect 13035 44152 14004 44180
rect 13035 44149 13047 44152
rect 12989 44143 13047 44149
rect 13998 44140 14004 44152
rect 14056 44140 14062 44192
rect 20070 44140 20076 44192
rect 20128 44140 20134 44192
rect 21008 44189 21036 44288
rect 20993 44183 21051 44189
rect 20993 44149 21005 44183
rect 21039 44180 21051 44183
rect 21174 44180 21180 44192
rect 21039 44152 21180 44180
rect 21039 44149 21051 44152
rect 20993 44143 21051 44149
rect 21174 44140 21180 44152
rect 21232 44140 21238 44192
rect 1104 44090 28888 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 28888 44090
rect 1104 44016 28888 44038
rect 7101 43979 7159 43985
rect 7101 43945 7113 43979
rect 7147 43976 7159 43979
rect 7466 43976 7472 43988
rect 7147 43948 7472 43976
rect 7147 43945 7159 43948
rect 7101 43939 7159 43945
rect 7466 43936 7472 43948
rect 7524 43936 7530 43988
rect 9585 43979 9643 43985
rect 9585 43945 9597 43979
rect 9631 43976 9643 43979
rect 11790 43976 11796 43988
rect 9631 43948 11796 43976
rect 9631 43945 9643 43948
rect 9585 43939 9643 43945
rect 11790 43936 11796 43948
rect 11848 43936 11854 43988
rect 11900 43948 12664 43976
rect 9858 43840 9864 43852
rect 8496 43812 9864 43840
rect 4433 43775 4491 43781
rect 4433 43741 4445 43775
rect 4479 43772 4491 43775
rect 4522 43772 4528 43784
rect 4479 43744 4528 43772
rect 4479 43741 4491 43744
rect 4433 43735 4491 43741
rect 4522 43732 4528 43744
rect 4580 43772 4586 43784
rect 7190 43772 7196 43784
rect 4580 43744 7196 43772
rect 4580 43732 4586 43744
rect 7190 43732 7196 43744
rect 7248 43772 7254 43784
rect 8496 43781 8524 43812
rect 9858 43800 9864 43812
rect 9916 43800 9922 43852
rect 11900 43784 11928 43948
rect 12526 43868 12532 43920
rect 12584 43868 12590 43920
rect 12437 43843 12495 43849
rect 12437 43809 12449 43843
rect 12483 43840 12495 43843
rect 12544 43840 12572 43868
rect 12483 43812 12572 43840
rect 12636 43840 12664 43948
rect 12894 43936 12900 43988
rect 12952 43936 12958 43988
rect 13354 43936 13360 43988
rect 13412 43936 13418 43988
rect 18046 43936 18052 43988
rect 18104 43976 18110 43988
rect 18141 43979 18199 43985
rect 18141 43976 18153 43979
rect 18104 43948 18153 43976
rect 18104 43936 18110 43948
rect 18141 43945 18153 43948
rect 18187 43945 18199 43979
rect 18141 43939 18199 43945
rect 20254 43936 20260 43988
rect 20312 43936 20318 43988
rect 20441 43979 20499 43985
rect 20441 43945 20453 43979
rect 20487 43976 20499 43979
rect 20622 43976 20628 43988
rect 20487 43948 20628 43976
rect 20487 43945 20499 43948
rect 20441 43939 20499 43945
rect 20622 43936 20628 43948
rect 20680 43936 20686 43988
rect 12710 43868 12716 43920
rect 12768 43908 12774 43920
rect 13170 43908 13176 43920
rect 12768 43880 13176 43908
rect 12768 43868 12774 43880
rect 13170 43868 13176 43880
rect 13228 43908 13234 43920
rect 13449 43911 13507 43917
rect 13449 43908 13461 43911
rect 13228 43880 13461 43908
rect 13228 43868 13234 43880
rect 13449 43877 13461 43880
rect 13495 43877 13507 43911
rect 14734 43908 14740 43920
rect 13449 43871 13507 43877
rect 13556 43880 14740 43908
rect 13556 43840 13584 43880
rect 14734 43868 14740 43880
rect 14792 43868 14798 43920
rect 17865 43911 17923 43917
rect 17865 43877 17877 43911
rect 17911 43908 17923 43911
rect 19334 43908 19340 43920
rect 17911 43880 19340 43908
rect 17911 43877 17923 43880
rect 17865 43871 17923 43877
rect 19334 43868 19340 43880
rect 19392 43868 19398 43920
rect 12636 43812 13584 43840
rect 12483 43809 12495 43812
rect 12437 43803 12495 43809
rect 13814 43800 13820 43852
rect 13872 43800 13878 43852
rect 14090 43800 14096 43852
rect 14148 43840 14154 43852
rect 14185 43843 14243 43849
rect 14185 43840 14197 43843
rect 14148 43812 14197 43840
rect 14148 43800 14154 43812
rect 14185 43809 14197 43812
rect 14231 43809 14243 43843
rect 14185 43803 14243 43809
rect 14366 43800 14372 43852
rect 14424 43840 14430 43852
rect 14461 43843 14519 43849
rect 14461 43840 14473 43843
rect 14424 43812 14473 43840
rect 14424 43800 14430 43812
rect 14461 43809 14473 43812
rect 14507 43809 14519 43843
rect 14461 43803 14519 43809
rect 15010 43800 15016 43852
rect 15068 43800 15074 43852
rect 20809 43843 20867 43849
rect 20809 43840 20821 43843
rect 17236 43812 19472 43840
rect 8481 43775 8539 43781
rect 8481 43772 8493 43775
rect 7248 43744 8493 43772
rect 7248 43732 7254 43744
rect 8481 43741 8493 43744
rect 8527 43741 8539 43775
rect 8481 43735 8539 43741
rect 9309 43775 9367 43781
rect 9309 43741 9321 43775
rect 9355 43741 9367 43775
rect 9309 43735 9367 43741
rect 9401 43775 9459 43781
rect 9401 43741 9413 43775
rect 9447 43772 9459 43775
rect 10962 43772 10968 43784
rect 9447 43744 10968 43772
rect 9447 43741 9459 43744
rect 9401 43735 9459 43741
rect 4706 43713 4712 43716
rect 4700 43704 4712 43713
rect 4667 43676 4712 43704
rect 4700 43667 4712 43676
rect 4706 43664 4712 43667
rect 4764 43664 4770 43716
rect 7834 43664 7840 43716
rect 7892 43704 7898 43716
rect 8214 43707 8272 43713
rect 8214 43704 8226 43707
rect 7892 43676 8226 43704
rect 7892 43664 7898 43676
rect 8214 43673 8226 43676
rect 8260 43673 8272 43707
rect 9324 43704 9352 43735
rect 10962 43732 10968 43744
rect 11020 43732 11026 43784
rect 11790 43732 11796 43784
rect 11848 43732 11854 43784
rect 11882 43732 11888 43784
rect 11940 43732 11946 43784
rect 11974 43732 11980 43784
rect 12032 43732 12038 43784
rect 12161 43775 12219 43781
rect 12161 43741 12173 43775
rect 12207 43772 12219 43775
rect 12250 43772 12256 43784
rect 12207 43744 12256 43772
rect 12207 43741 12219 43744
rect 12161 43735 12219 43741
rect 12250 43732 12256 43744
rect 12308 43732 12314 43784
rect 12529 43775 12587 43781
rect 12529 43741 12541 43775
rect 12575 43741 12587 43775
rect 12529 43735 12587 43741
rect 12713 43775 12771 43781
rect 12713 43741 12725 43775
rect 12759 43772 12771 43775
rect 13538 43772 13544 43784
rect 12759 43744 13544 43772
rect 12759 43741 12771 43744
rect 12713 43735 12771 43741
rect 9950 43704 9956 43716
rect 9324 43676 9956 43704
rect 8214 43667 8272 43673
rect 9950 43664 9956 43676
rect 10008 43664 10014 43716
rect 10128 43707 10186 43713
rect 10128 43673 10140 43707
rect 10174 43704 10186 43707
rect 11517 43707 11575 43713
rect 11517 43704 11529 43707
rect 10174 43676 11529 43704
rect 10174 43673 10186 43676
rect 10128 43667 10186 43673
rect 11517 43673 11529 43676
rect 11563 43673 11575 43707
rect 11808 43704 11836 43732
rect 12544 43704 12572 43735
rect 13538 43732 13544 43744
rect 13596 43772 13602 43784
rect 14384 43772 14412 43800
rect 13596 43744 14412 43772
rect 14553 43775 14611 43781
rect 13596 43732 13602 43744
rect 14553 43741 14565 43775
rect 14599 43772 14611 43775
rect 15562 43772 15568 43784
rect 14599 43744 15568 43772
rect 14599 43741 14611 43744
rect 14553 43735 14611 43741
rect 15562 43732 15568 43744
rect 15620 43732 15626 43784
rect 16666 43732 16672 43784
rect 16724 43732 16730 43784
rect 16758 43732 16764 43784
rect 16816 43732 16822 43784
rect 17126 43732 17132 43784
rect 17184 43781 17190 43784
rect 17184 43772 17192 43781
rect 17236 43772 17264 43812
rect 17589 43775 17647 43781
rect 17589 43772 17601 43775
rect 17184 43744 17264 43772
rect 17328 43744 17601 43772
rect 17184 43735 17192 43744
rect 17184 43732 17190 43735
rect 11808 43676 12572 43704
rect 15280 43707 15338 43713
rect 11517 43667 11575 43673
rect 15280 43673 15292 43707
rect 15326 43704 15338 43707
rect 15838 43704 15844 43716
rect 15326 43676 15844 43704
rect 15326 43673 15338 43676
rect 15280 43667 15338 43673
rect 15838 43664 15844 43676
rect 15896 43664 15902 43716
rect 16850 43704 16856 43716
rect 16408 43676 16856 43704
rect 16408 43648 16436 43676
rect 16850 43664 16856 43676
rect 16908 43664 16914 43716
rect 16942 43664 16948 43716
rect 17000 43664 17006 43716
rect 17037 43707 17095 43713
rect 17037 43673 17049 43707
rect 17083 43673 17095 43707
rect 17037 43667 17095 43673
rect 5813 43639 5871 43645
rect 5813 43605 5825 43639
rect 5859 43636 5871 43639
rect 6454 43636 6460 43648
rect 5859 43608 6460 43636
rect 5859 43605 5871 43608
rect 5813 43599 5871 43605
rect 6454 43596 6460 43608
rect 6512 43596 6518 43648
rect 11241 43639 11299 43645
rect 11241 43605 11253 43639
rect 11287 43636 11299 43639
rect 11606 43636 11612 43648
rect 11287 43608 11612 43636
rect 11287 43605 11299 43608
rect 11241 43599 11299 43605
rect 11606 43596 11612 43608
rect 11664 43596 11670 43648
rect 16390 43596 16396 43648
rect 16448 43596 16454 43648
rect 16482 43596 16488 43648
rect 16540 43636 16546 43648
rect 17052 43636 17080 43667
rect 17218 43636 17224 43648
rect 16540 43608 17224 43636
rect 16540 43596 16546 43608
rect 17218 43596 17224 43608
rect 17276 43596 17282 43648
rect 17328 43645 17356 43744
rect 17589 43741 17601 43744
rect 17635 43741 17647 43775
rect 17589 43735 17647 43741
rect 17678 43732 17684 43784
rect 17736 43732 17742 43784
rect 18785 43775 18843 43781
rect 18785 43741 18797 43775
rect 18831 43772 18843 43775
rect 19337 43775 19395 43781
rect 19337 43772 19349 43775
rect 18831 43744 19349 43772
rect 18831 43741 18843 43744
rect 18785 43735 18843 43741
rect 19337 43741 19349 43744
rect 19383 43741 19395 43775
rect 19337 43735 19395 43741
rect 17862 43664 17868 43716
rect 17920 43664 17926 43716
rect 19444 43704 19472 43812
rect 19536 43812 20821 43840
rect 19536 43781 19564 43812
rect 20809 43809 20821 43812
rect 20855 43809 20867 43843
rect 20809 43803 20867 43809
rect 19521 43775 19579 43781
rect 19521 43741 19533 43775
rect 19567 43741 19579 43775
rect 19521 43735 19579 43741
rect 19702 43732 19708 43784
rect 19760 43732 19766 43784
rect 19797 43775 19855 43781
rect 19797 43741 19809 43775
rect 19843 43741 19855 43775
rect 19797 43735 19855 43741
rect 19812 43704 19840 43735
rect 20622 43732 20628 43784
rect 20680 43772 20686 43784
rect 20717 43775 20775 43781
rect 20717 43772 20729 43775
rect 20680 43744 20729 43772
rect 20680 43732 20686 43744
rect 20717 43741 20729 43744
rect 20763 43741 20775 43775
rect 20717 43735 20775 43741
rect 20901 43775 20959 43781
rect 20901 43741 20913 43775
rect 20947 43772 20959 43775
rect 20947 43744 21220 43772
rect 20947 43741 20959 43744
rect 20901 43735 20959 43741
rect 20070 43704 20076 43716
rect 19444 43676 20076 43704
rect 20070 43664 20076 43676
rect 20128 43664 20134 43716
rect 21192 43648 21220 43744
rect 17313 43639 17371 43645
rect 17313 43605 17325 43639
rect 17359 43605 17371 43639
rect 17313 43599 17371 43605
rect 19242 43596 19248 43648
rect 19300 43636 19306 43648
rect 20273 43639 20331 43645
rect 20273 43636 20285 43639
rect 19300 43608 20285 43636
rect 19300 43596 19306 43608
rect 20273 43605 20285 43608
rect 20319 43605 20331 43639
rect 20273 43599 20331 43605
rect 21174 43596 21180 43648
rect 21232 43596 21238 43648
rect 1104 43546 28888 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 28888 43546
rect 1104 43472 28888 43494
rect 11057 43435 11115 43441
rect 11057 43401 11069 43435
rect 11103 43432 11115 43435
rect 11974 43432 11980 43444
rect 11103 43404 11980 43432
rect 11103 43401 11115 43404
rect 11057 43395 11115 43401
rect 11974 43392 11980 43404
rect 12032 43392 12038 43444
rect 13170 43392 13176 43444
rect 13228 43392 13234 43444
rect 15838 43392 15844 43444
rect 15896 43392 15902 43444
rect 16758 43392 16764 43444
rect 16816 43392 16822 43444
rect 18414 43392 18420 43444
rect 18472 43432 18478 43444
rect 20254 43432 20260 43444
rect 18472 43404 20260 43432
rect 18472 43392 18478 43404
rect 20254 43392 20260 43404
rect 20312 43432 20318 43444
rect 20533 43435 20591 43441
rect 20533 43432 20545 43435
rect 20312 43404 20545 43432
rect 20312 43392 20318 43404
rect 20533 43401 20545 43404
rect 20579 43401 20591 43435
rect 20533 43395 20591 43401
rect 10413 43367 10471 43373
rect 10413 43333 10425 43367
rect 10459 43364 10471 43367
rect 11882 43364 11888 43376
rect 10459 43336 11888 43364
rect 10459 43333 10471 43336
rect 10413 43327 10471 43333
rect 11882 43324 11888 43336
rect 11940 43324 11946 43376
rect 13357 43367 13415 43373
rect 13357 43333 13369 43367
rect 13403 43364 13415 43367
rect 13906 43364 13912 43376
rect 13403 43336 13912 43364
rect 13403 43333 13415 43336
rect 13357 43327 13415 43333
rect 13906 43324 13912 43336
rect 13964 43324 13970 43376
rect 18432 43364 18460 43392
rect 16960 43336 18460 43364
rect 6454 43256 6460 43308
rect 6512 43256 6518 43308
rect 10042 43256 10048 43308
rect 10100 43296 10106 43308
rect 10781 43299 10839 43305
rect 10781 43296 10793 43299
rect 10100 43268 10793 43296
rect 10100 43256 10106 43268
rect 10781 43265 10793 43268
rect 10827 43265 10839 43299
rect 10781 43259 10839 43265
rect 10873 43299 10931 43305
rect 10873 43265 10885 43299
rect 10919 43296 10931 43299
rect 11054 43296 11060 43308
rect 10919 43268 11060 43296
rect 10919 43265 10931 43268
rect 10873 43259 10931 43265
rect 11054 43256 11060 43268
rect 11112 43256 11118 43308
rect 11606 43256 11612 43308
rect 11664 43296 11670 43308
rect 11664 43268 12434 43296
rect 11664 43256 11670 43268
rect 12406 43228 12434 43268
rect 12526 43256 12532 43308
rect 12584 43256 12590 43308
rect 13538 43256 13544 43308
rect 13596 43256 13602 43308
rect 13998 43256 14004 43308
rect 14056 43256 14062 43308
rect 16960 43305 16988 43336
rect 16945 43299 17003 43305
rect 16945 43265 16957 43299
rect 16991 43265 17003 43299
rect 16945 43259 17003 43265
rect 17034 43256 17040 43308
rect 17092 43256 17098 43308
rect 17218 43256 17224 43308
rect 17276 43296 17282 43308
rect 17696 43305 17724 43336
rect 17313 43299 17371 43305
rect 17313 43296 17325 43299
rect 17276 43268 17325 43296
rect 17276 43256 17282 43268
rect 17313 43265 17325 43268
rect 17359 43265 17371 43299
rect 17313 43259 17371 43265
rect 17681 43299 17739 43305
rect 17681 43265 17693 43299
rect 17727 43265 17739 43299
rect 17681 43259 17739 43265
rect 17773 43299 17831 43305
rect 17773 43265 17785 43299
rect 17819 43296 17831 43299
rect 17954 43296 17960 43308
rect 17819 43268 17960 43296
rect 17819 43265 17831 43268
rect 17773 43259 17831 43265
rect 17954 43256 17960 43268
rect 18012 43256 18018 43308
rect 18230 43256 18236 43308
rect 18288 43256 18294 43308
rect 18500 43299 18558 43305
rect 18500 43265 18512 43299
rect 18546 43296 18558 43299
rect 19334 43296 19340 43308
rect 18546 43268 19340 43296
rect 18546 43265 18558 43268
rect 18500 43259 18558 43265
rect 19334 43256 19340 43268
rect 19392 43256 19398 43308
rect 12618 43228 12624 43240
rect 12406 43200 12624 43228
rect 12618 43188 12624 43200
rect 12676 43188 12682 43240
rect 14090 43188 14096 43240
rect 14148 43188 14154 43240
rect 15194 43188 15200 43240
rect 15252 43188 15258 43240
rect 19889 43231 19947 43237
rect 19889 43228 19901 43231
rect 19628 43200 19901 43228
rect 11974 43120 11980 43172
rect 12032 43160 12038 43172
rect 14369 43163 14427 43169
rect 12032 43132 12664 43160
rect 12032 43120 12038 43132
rect 5810 43052 5816 43104
rect 5868 43092 5874 43104
rect 6822 43092 6828 43104
rect 5868 43064 6828 43092
rect 5868 43052 5874 43064
rect 6822 43052 6828 43064
rect 6880 43092 6886 43104
rect 7101 43095 7159 43101
rect 7101 43092 7113 43095
rect 6880 43064 7113 43092
rect 6880 43052 6886 43064
rect 7101 43061 7113 43064
rect 7147 43061 7159 43095
rect 7101 43055 7159 43061
rect 11790 43052 11796 43104
rect 11848 43092 11854 43104
rect 12253 43095 12311 43101
rect 12253 43092 12265 43095
rect 11848 43064 12265 43092
rect 11848 43052 11854 43064
rect 12253 43061 12265 43064
rect 12299 43092 12311 43095
rect 12434 43092 12440 43104
rect 12299 43064 12440 43092
rect 12299 43061 12311 43064
rect 12253 43055 12311 43061
rect 12434 43052 12440 43064
rect 12492 43052 12498 43104
rect 12636 43101 12664 43132
rect 14369 43129 14381 43163
rect 14415 43160 14427 43163
rect 14642 43160 14648 43172
rect 14415 43132 14648 43160
rect 14415 43129 14427 43132
rect 14369 43123 14427 43129
rect 14642 43120 14648 43132
rect 14700 43120 14706 43172
rect 17126 43120 17132 43172
rect 17184 43160 17190 43172
rect 19628 43169 19656 43200
rect 19889 43197 19901 43200
rect 19935 43197 19947 43231
rect 19889 43191 19947 43197
rect 17221 43163 17279 43169
rect 17221 43160 17233 43163
rect 17184 43132 17233 43160
rect 17184 43120 17190 43132
rect 17221 43129 17233 43132
rect 17267 43129 17279 43163
rect 17221 43123 17279 43129
rect 19613 43163 19671 43169
rect 19613 43129 19625 43163
rect 19659 43129 19671 43163
rect 19613 43123 19671 43129
rect 12621 43095 12679 43101
rect 12621 43061 12633 43095
rect 12667 43092 12679 43095
rect 17034 43092 17040 43104
rect 12667 43064 17040 43092
rect 12667 43061 12679 43064
rect 12621 43055 12679 43061
rect 17034 43052 17040 43064
rect 17092 43052 17098 43104
rect 17957 43095 18015 43101
rect 17957 43061 17969 43095
rect 18003 43092 18015 43095
rect 19702 43092 19708 43104
rect 18003 43064 19708 43092
rect 18003 43061 18015 43064
rect 17957 43055 18015 43061
rect 19702 43052 19708 43064
rect 19760 43052 19766 43104
rect 1104 43002 28888 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 28888 43002
rect 1104 42928 28888 42950
rect 11698 42848 11704 42900
rect 11756 42848 11762 42900
rect 12529 42891 12587 42897
rect 12529 42888 12541 42891
rect 12406 42860 12541 42888
rect 9950 42780 9956 42832
rect 10008 42820 10014 42832
rect 12406 42820 12434 42860
rect 12529 42857 12541 42860
rect 12575 42857 12587 42891
rect 12529 42851 12587 42857
rect 16669 42891 16727 42897
rect 16669 42857 16681 42891
rect 16715 42888 16727 42891
rect 16942 42888 16948 42900
rect 16715 42860 16948 42888
rect 16715 42857 16727 42860
rect 16669 42851 16727 42857
rect 16942 42848 16948 42860
rect 17000 42848 17006 42900
rect 10008 42792 12434 42820
rect 10008 42780 10014 42792
rect 17954 42780 17960 42832
rect 18012 42820 18018 42832
rect 18877 42823 18935 42829
rect 18012 42792 18552 42820
rect 18012 42780 18018 42792
rect 10962 42712 10968 42764
rect 11020 42712 11026 42764
rect 11330 42712 11336 42764
rect 11388 42752 11394 42764
rect 12066 42752 12072 42764
rect 11388 42724 12072 42752
rect 11388 42712 11394 42724
rect 12066 42712 12072 42724
rect 12124 42752 12130 42764
rect 14277 42755 14335 42761
rect 12124 42724 12664 42752
rect 12124 42712 12130 42724
rect 4706 42644 4712 42696
rect 4764 42684 4770 42696
rect 5077 42687 5135 42693
rect 5077 42684 5089 42687
rect 4764 42656 5089 42684
rect 4764 42644 4770 42656
rect 5077 42653 5089 42656
rect 5123 42653 5135 42687
rect 5077 42647 5135 42653
rect 11149 42687 11207 42693
rect 11149 42653 11161 42687
rect 11195 42684 11207 42687
rect 11790 42684 11796 42696
rect 11195 42656 11796 42684
rect 11195 42653 11207 42656
rect 11149 42647 11207 42653
rect 11790 42644 11796 42656
rect 11848 42644 11854 42696
rect 11974 42693 11980 42696
rect 11931 42687 11980 42693
rect 11931 42653 11943 42687
rect 11977 42653 11980 42687
rect 11931 42647 11980 42653
rect 11974 42644 11980 42647
rect 12032 42644 12038 42696
rect 12434 42644 12440 42696
rect 12492 42644 12498 42696
rect 12636 42693 12664 42724
rect 14277 42721 14289 42755
rect 14323 42752 14335 42755
rect 14921 42755 14979 42761
rect 14921 42752 14933 42755
rect 14323 42724 14933 42752
rect 14323 42721 14335 42724
rect 14277 42715 14335 42721
rect 14921 42721 14933 42724
rect 14967 42721 14979 42755
rect 14921 42715 14979 42721
rect 15105 42755 15163 42761
rect 15105 42721 15117 42755
rect 15151 42752 15163 42755
rect 15194 42752 15200 42764
rect 15151 42724 15200 42752
rect 15151 42721 15163 42724
rect 15105 42715 15163 42721
rect 15194 42712 15200 42724
rect 15252 42712 15258 42764
rect 18414 42712 18420 42764
rect 18472 42712 18478 42764
rect 18524 42761 18552 42792
rect 18877 42789 18889 42823
rect 18923 42820 18935 42823
rect 18923 42792 19932 42820
rect 18923 42789 18935 42792
rect 18877 42783 18935 42789
rect 18509 42755 18567 42761
rect 18509 42721 18521 42755
rect 18555 42752 18567 42755
rect 19242 42752 19248 42764
rect 18555 42724 19248 42752
rect 18555 42721 18567 42724
rect 18509 42715 18567 42721
rect 19242 42712 19248 42724
rect 19300 42712 19306 42764
rect 19334 42712 19340 42764
rect 19392 42712 19398 42764
rect 19904 42761 19932 42792
rect 19889 42755 19947 42761
rect 19889 42721 19901 42755
rect 19935 42721 19947 42755
rect 19889 42715 19947 42721
rect 12621 42687 12679 42693
rect 12621 42653 12633 42687
rect 12667 42684 12679 42687
rect 13538 42684 13544 42696
rect 12667 42656 13544 42684
rect 12667 42653 12679 42656
rect 12621 42647 12679 42653
rect 13538 42644 13544 42656
rect 13596 42644 13602 42696
rect 14090 42644 14096 42696
rect 14148 42684 14154 42696
rect 14185 42687 14243 42693
rect 14185 42684 14197 42687
rect 14148 42656 14197 42684
rect 14148 42644 14154 42656
rect 14185 42653 14197 42656
rect 14231 42653 14243 42687
rect 14185 42647 14243 42653
rect 14369 42687 14427 42693
rect 14369 42653 14381 42687
rect 14415 42653 14427 42687
rect 14369 42647 14427 42653
rect 5344 42619 5402 42625
rect 5344 42585 5356 42619
rect 5390 42616 5402 42619
rect 5442 42616 5448 42628
rect 5390 42588 5448 42616
rect 5390 42585 5402 42588
rect 5344 42579 5402 42585
rect 5442 42576 5448 42588
rect 5500 42576 5506 42628
rect 11330 42576 11336 42628
rect 11388 42576 11394 42628
rect 6454 42508 6460 42560
rect 6512 42508 6518 42560
rect 14200 42548 14228 42647
rect 14384 42616 14412 42647
rect 14642 42644 14648 42696
rect 14700 42644 14706 42696
rect 15010 42644 15016 42696
rect 15068 42684 15074 42696
rect 15068 42656 15700 42684
rect 15068 42644 15074 42656
rect 15562 42616 15568 42628
rect 14384 42588 15568 42616
rect 15562 42576 15568 42588
rect 15620 42576 15626 42628
rect 14734 42548 14740 42560
rect 14200 42520 14740 42548
rect 14734 42508 14740 42520
rect 14792 42508 14798 42560
rect 15473 42551 15531 42557
rect 15473 42517 15485 42551
rect 15519 42548 15531 42551
rect 15672 42548 15700 42656
rect 16114 42644 16120 42696
rect 16172 42644 16178 42696
rect 16485 42687 16543 42693
rect 16485 42653 16497 42687
rect 16531 42684 16543 42687
rect 18432 42684 18460 42712
rect 16531 42656 18460 42684
rect 18693 42687 18751 42693
rect 16531 42653 16543 42656
rect 16485 42647 16543 42653
rect 18693 42653 18705 42687
rect 18739 42684 18751 42687
rect 19426 42684 19432 42696
rect 18739 42656 19432 42684
rect 18739 42653 18751 42656
rect 18693 42647 18751 42653
rect 19426 42644 19432 42656
rect 19484 42644 19490 42696
rect 16298 42576 16304 42628
rect 16356 42576 16362 42628
rect 16393 42619 16451 42625
rect 16393 42585 16405 42619
rect 16439 42616 16451 42619
rect 17034 42616 17040 42628
rect 16439 42588 17040 42616
rect 16439 42585 16451 42588
rect 16393 42579 16451 42585
rect 17034 42576 17040 42588
rect 17092 42576 17098 42628
rect 16482 42548 16488 42560
rect 15519 42520 16488 42548
rect 15519 42517 15531 42520
rect 15473 42511 15531 42517
rect 16482 42508 16488 42520
rect 16540 42548 16546 42560
rect 17862 42548 17868 42560
rect 16540 42520 17868 42548
rect 16540 42508 16546 42520
rect 17862 42508 17868 42520
rect 17920 42548 17926 42560
rect 17957 42551 18015 42557
rect 17957 42548 17969 42551
rect 17920 42520 17969 42548
rect 17920 42508 17926 42520
rect 17957 42517 17969 42520
rect 18003 42517 18015 42551
rect 17957 42511 18015 42517
rect 1104 42458 28888 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 28888 42458
rect 1104 42384 28888 42406
rect 5442 42304 5448 42356
rect 5500 42304 5506 42356
rect 19426 42304 19432 42356
rect 19484 42304 19490 42356
rect 19702 42276 19708 42288
rect 19352 42248 19708 42276
rect 5626 42168 5632 42220
rect 5684 42168 5690 42220
rect 5810 42168 5816 42220
rect 5868 42168 5874 42220
rect 6454 42168 6460 42220
rect 6512 42168 6518 42220
rect 19352 42217 19380 42248
rect 19702 42236 19708 42248
rect 19760 42236 19766 42288
rect 19337 42211 19395 42217
rect 19337 42177 19349 42211
rect 19383 42177 19395 42211
rect 19337 42171 19395 42177
rect 19521 42211 19579 42217
rect 19521 42177 19533 42211
rect 19567 42208 19579 42211
rect 19567 42180 19932 42208
rect 19567 42177 19579 42180
rect 19521 42171 19579 42177
rect 7098 41964 7104 42016
rect 7156 41964 7162 42016
rect 19904 42013 19932 42180
rect 19889 42007 19947 42013
rect 19889 41973 19901 42007
rect 19935 42004 19947 42007
rect 20162 42004 20168 42016
rect 19935 41976 20168 42004
rect 19935 41973 19947 41976
rect 19889 41967 19947 41973
rect 20162 41964 20168 41976
rect 20220 42004 20226 42016
rect 21174 42004 21180 42016
rect 20220 41976 21180 42004
rect 20220 41964 20226 41976
rect 21174 41964 21180 41976
rect 21232 41964 21238 42016
rect 1104 41914 28888 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 28888 41914
rect 1104 41840 28888 41862
rect 5997 41667 6055 41673
rect 5997 41633 6009 41667
rect 6043 41664 6055 41667
rect 7098 41664 7104 41676
rect 6043 41636 7104 41664
rect 6043 41633 6055 41636
rect 5997 41627 6055 41633
rect 7098 41624 7104 41636
rect 7156 41624 7162 41676
rect 5626 41556 5632 41608
rect 5684 41596 5690 41608
rect 5813 41599 5871 41605
rect 5813 41596 5825 41599
rect 5684 41568 5825 41596
rect 5684 41556 5690 41568
rect 5813 41565 5825 41568
rect 5859 41565 5871 41599
rect 5813 41559 5871 41565
rect 12618 41556 12624 41608
rect 12676 41596 12682 41608
rect 13541 41599 13599 41605
rect 13541 41596 13553 41599
rect 12676 41568 13553 41596
rect 12676 41556 12682 41568
rect 13541 41565 13553 41568
rect 13587 41565 13599 41599
rect 13541 41559 13599 41565
rect 5534 41420 5540 41472
rect 5592 41460 5598 41472
rect 5629 41463 5687 41469
rect 5629 41460 5641 41463
rect 5592 41432 5641 41460
rect 5592 41420 5598 41432
rect 5629 41429 5641 41432
rect 5675 41429 5687 41463
rect 5629 41423 5687 41429
rect 13633 41463 13691 41469
rect 13633 41429 13645 41463
rect 13679 41460 13691 41463
rect 16022 41460 16028 41472
rect 13679 41432 16028 41460
rect 13679 41429 13691 41432
rect 13633 41423 13691 41429
rect 16022 41420 16028 41432
rect 16080 41420 16086 41472
rect 1104 41370 28888 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 28888 41370
rect 1104 41296 28888 41318
rect 6822 41216 6828 41268
rect 6880 41256 6886 41268
rect 7561 41259 7619 41265
rect 7561 41256 7573 41259
rect 6880 41228 7573 41256
rect 6880 41216 6886 41228
rect 7561 41225 7573 41228
rect 7607 41225 7619 41259
rect 7561 41219 7619 41225
rect 5442 41188 5448 41200
rect 4724 41160 5448 41188
rect 4724 41132 4752 41160
rect 5442 41148 5448 41160
rect 5500 41148 5506 41200
rect 6638 41148 6644 41200
rect 6696 41188 6702 41200
rect 6696 41160 6914 41188
rect 6696 41148 6702 41160
rect 4706 41080 4712 41132
rect 4764 41080 4770 41132
rect 4976 41123 5034 41129
rect 4976 41089 4988 41123
rect 5022 41120 5034 41123
rect 5534 41120 5540 41132
rect 5022 41092 5540 41120
rect 5022 41089 5034 41092
rect 4976 41083 5034 41089
rect 5534 41080 5540 41092
rect 5592 41080 5598 41132
rect 6886 41120 6914 41160
rect 7190 41148 7196 41200
rect 7248 41188 7254 41200
rect 7377 41191 7435 41197
rect 7377 41188 7389 41191
rect 7248 41160 7389 41188
rect 7248 41148 7254 41160
rect 7377 41157 7389 41160
rect 7423 41157 7435 41191
rect 7377 41151 7435 41157
rect 7101 41123 7159 41129
rect 7101 41120 7113 41123
rect 6886 41092 7113 41120
rect 7101 41089 7113 41092
rect 7147 41120 7159 41123
rect 7653 41123 7711 41129
rect 7653 41120 7665 41123
rect 7147 41092 7665 41120
rect 7147 41089 7159 41092
rect 7101 41083 7159 41089
rect 7653 41089 7665 41092
rect 7699 41089 7711 41123
rect 7653 41083 7711 41089
rect 7745 41123 7803 41129
rect 7745 41089 7757 41123
rect 7791 41120 7803 41123
rect 7926 41120 7932 41132
rect 7791 41092 7932 41120
rect 7791 41089 7803 41092
rect 7745 41083 7803 41089
rect 7926 41080 7932 41092
rect 7984 41080 7990 41132
rect 6457 41055 6515 41061
rect 6457 41021 6469 41055
rect 6503 41021 6515 41055
rect 6457 41015 6515 41021
rect 6089 40987 6147 40993
rect 6089 40953 6101 40987
rect 6135 40984 6147 40987
rect 6472 40984 6500 41015
rect 6135 40956 6500 40984
rect 6135 40953 6147 40956
rect 6089 40947 6147 40953
rect 7466 40876 7472 40928
rect 7524 40916 7530 40928
rect 7929 40919 7987 40925
rect 7929 40916 7941 40919
rect 7524 40888 7941 40916
rect 7524 40876 7530 40888
rect 7929 40885 7941 40888
rect 7975 40885 7987 40919
rect 7929 40879 7987 40885
rect 1104 40826 28888 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 28888 40826
rect 1104 40752 28888 40774
rect 6822 40672 6828 40724
rect 6880 40672 6886 40724
rect 7742 40672 7748 40724
rect 7800 40712 7806 40724
rect 8113 40715 8171 40721
rect 8113 40712 8125 40715
rect 7800 40684 8125 40712
rect 7800 40672 7806 40684
rect 8113 40681 8125 40684
rect 8159 40712 8171 40715
rect 8570 40712 8576 40724
rect 8159 40684 8576 40712
rect 8159 40681 8171 40684
rect 8113 40675 8171 40681
rect 8570 40672 8576 40684
rect 8628 40672 8634 40724
rect 9490 40672 9496 40724
rect 9548 40712 9554 40724
rect 10686 40712 10692 40724
rect 9548 40684 10692 40712
rect 9548 40672 9554 40684
rect 10686 40672 10692 40684
rect 10744 40672 10750 40724
rect 16209 40715 16267 40721
rect 16209 40681 16221 40715
rect 16255 40712 16267 40715
rect 16298 40712 16304 40724
rect 16255 40684 16304 40712
rect 16255 40681 16267 40684
rect 16209 40675 16267 40681
rect 16298 40672 16304 40684
rect 16356 40672 16362 40724
rect 8297 40647 8355 40653
rect 8297 40613 8309 40647
rect 8343 40644 8355 40647
rect 10870 40644 10876 40656
rect 8343 40616 10876 40644
rect 8343 40613 8355 40616
rect 8297 40607 8355 40613
rect 10870 40604 10876 40616
rect 10928 40604 10934 40656
rect 6825 40579 6883 40585
rect 6825 40545 6837 40579
rect 6871 40576 6883 40579
rect 7650 40576 7656 40588
rect 6871 40548 7656 40576
rect 6871 40545 6883 40548
rect 6825 40539 6883 40545
rect 7650 40536 7656 40548
rect 7708 40536 7714 40588
rect 7834 40536 7840 40588
rect 7892 40536 7898 40588
rect 7926 40536 7932 40588
rect 7984 40536 7990 40588
rect 5626 40468 5632 40520
rect 5684 40508 5690 40520
rect 6089 40511 6147 40517
rect 6089 40508 6101 40511
rect 5684 40480 6101 40508
rect 5684 40468 5690 40480
rect 6089 40477 6101 40480
rect 6135 40477 6147 40511
rect 6089 40471 6147 40477
rect 6273 40511 6331 40517
rect 6273 40477 6285 40511
rect 6319 40508 6331 40511
rect 6638 40508 6644 40520
rect 6319 40480 6644 40508
rect 6319 40477 6331 40480
rect 6273 40471 6331 40477
rect 6104 40440 6132 40471
rect 6638 40468 6644 40480
rect 6696 40468 6702 40520
rect 6917 40511 6975 40517
rect 6917 40477 6929 40511
rect 6963 40508 6975 40511
rect 7098 40508 7104 40520
rect 6963 40480 7104 40508
rect 6963 40477 6975 40480
rect 6917 40471 6975 40477
rect 7098 40468 7104 40480
rect 7156 40468 7162 40520
rect 7852 40508 7880 40536
rect 8113 40511 8171 40517
rect 8113 40508 8125 40511
rect 7852 40480 8125 40508
rect 8113 40477 8125 40480
rect 8159 40477 8171 40511
rect 8113 40471 8171 40477
rect 10137 40511 10195 40517
rect 10137 40477 10149 40511
rect 10183 40508 10195 40511
rect 10962 40508 10968 40520
rect 10183 40480 10968 40508
rect 10183 40477 10195 40480
rect 10137 40471 10195 40477
rect 10962 40468 10968 40480
rect 11020 40468 11026 40520
rect 16022 40468 16028 40520
rect 16080 40468 16086 40520
rect 7282 40440 7288 40452
rect 6104 40412 7288 40440
rect 7282 40400 7288 40412
rect 7340 40400 7346 40452
rect 7837 40443 7895 40449
rect 7837 40409 7849 40443
rect 7883 40409 7895 40443
rect 7837 40403 7895 40409
rect 5902 40332 5908 40384
rect 5960 40332 5966 40384
rect 7101 40375 7159 40381
rect 7101 40341 7113 40375
rect 7147 40372 7159 40375
rect 7852 40372 7880 40403
rect 15838 40400 15844 40452
rect 15896 40400 15902 40452
rect 7147 40344 7880 40372
rect 7147 40341 7159 40344
rect 7101 40335 7159 40341
rect 1104 40282 28888 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 28888 40282
rect 1104 40208 28888 40230
rect 7650 40128 7656 40180
rect 7708 40128 7714 40180
rect 7834 40128 7840 40180
rect 7892 40168 7898 40180
rect 9309 40171 9367 40177
rect 9309 40168 9321 40171
rect 7892 40140 9321 40168
rect 7892 40128 7898 40140
rect 9309 40137 9321 40140
rect 9355 40137 9367 40171
rect 9309 40131 9367 40137
rect 10962 40128 10968 40180
rect 11020 40128 11026 40180
rect 11606 40128 11612 40180
rect 11664 40128 11670 40180
rect 16025 40171 16083 40177
rect 16025 40137 16037 40171
rect 16071 40168 16083 40171
rect 16206 40168 16212 40180
rect 16071 40140 16212 40168
rect 16071 40137 16083 40140
rect 16025 40131 16083 40137
rect 16206 40128 16212 40140
rect 16264 40168 16270 40180
rect 16666 40168 16672 40180
rect 16264 40140 16672 40168
rect 16264 40128 16270 40140
rect 16666 40128 16672 40140
rect 16724 40128 16730 40180
rect 8128 40072 8340 40100
rect 7929 40035 7987 40041
rect 7929 40001 7941 40035
rect 7975 40032 7987 40035
rect 8018 40032 8024 40044
rect 7975 40004 8024 40032
rect 7975 40001 7987 40004
rect 7929 39995 7987 40001
rect 8018 39992 8024 40004
rect 8076 40032 8082 40044
rect 8128 40032 8156 40072
rect 8202 40041 8208 40044
rect 8076 40004 8156 40032
rect 8076 39992 8082 40004
rect 8196 39995 8208 40041
rect 8202 39992 8208 39995
rect 8260 39992 8266 40044
rect 8312 40032 8340 40072
rect 9585 40035 9643 40041
rect 9585 40032 9597 40035
rect 8312 40004 9597 40032
rect 9585 40001 9597 40004
rect 9631 40001 9643 40035
rect 9585 39995 9643 40001
rect 9674 39992 9680 40044
rect 9732 40032 9738 40044
rect 9841 40035 9899 40041
rect 9841 40032 9853 40035
rect 9732 40004 9853 40032
rect 9732 39992 9738 40004
rect 9841 40001 9853 40004
rect 9887 40001 9899 40035
rect 9841 39995 9899 40001
rect 11238 39992 11244 40044
rect 11296 40032 11302 40044
rect 11977 40035 12035 40041
rect 11977 40032 11989 40035
rect 11296 40004 11989 40032
rect 11296 39992 11302 40004
rect 11977 40001 11989 40004
rect 12023 40001 12035 40035
rect 11977 39995 12035 40001
rect 14552 40035 14610 40041
rect 14552 40001 14564 40035
rect 14598 40001 14610 40035
rect 14552 39995 14610 40001
rect 14645 40035 14703 40041
rect 14645 40001 14657 40035
rect 14691 40032 14703 40035
rect 15286 40032 15292 40044
rect 14691 40004 15292 40032
rect 14691 40001 14703 40004
rect 14645 39995 14703 40001
rect 7006 39924 7012 39976
rect 7064 39924 7070 39976
rect 11422 39924 11428 39976
rect 11480 39964 11486 39976
rect 11793 39967 11851 39973
rect 11793 39964 11805 39967
rect 11480 39936 11805 39964
rect 11480 39924 11486 39936
rect 11793 39933 11805 39936
rect 11839 39933 11851 39967
rect 11793 39927 11851 39933
rect 11885 39967 11943 39973
rect 11885 39933 11897 39967
rect 11931 39933 11943 39967
rect 11885 39927 11943 39933
rect 12069 39967 12127 39973
rect 12069 39933 12081 39967
rect 12115 39964 12127 39967
rect 13170 39964 13176 39976
rect 12115 39936 13176 39964
rect 12115 39933 12127 39936
rect 12069 39927 12127 39933
rect 11146 39856 11152 39908
rect 11204 39896 11210 39908
rect 11900 39896 11928 39927
rect 13170 39924 13176 39936
rect 13228 39924 13234 39976
rect 14568 39964 14596 39995
rect 15286 39992 15292 40004
rect 15344 39992 15350 40044
rect 15562 39992 15568 40044
rect 15620 39992 15626 40044
rect 15194 39964 15200 39976
rect 14568 39936 15200 39964
rect 15194 39924 15200 39936
rect 15252 39924 15258 39976
rect 17862 39924 17868 39976
rect 17920 39964 17926 39976
rect 18233 39967 18291 39973
rect 18233 39964 18245 39967
rect 17920 39936 18245 39964
rect 17920 39924 17926 39936
rect 18233 39933 18245 39936
rect 18279 39933 18291 39967
rect 18233 39927 18291 39933
rect 11204 39868 11928 39896
rect 11204 39856 11210 39868
rect 15746 39856 15752 39908
rect 15804 39896 15810 39908
rect 15841 39899 15899 39905
rect 15841 39896 15853 39899
rect 15804 39868 15853 39896
rect 15804 39856 15810 39868
rect 15841 39865 15853 39868
rect 15887 39865 15899 39899
rect 15841 39859 15899 39865
rect 14461 39831 14519 39837
rect 14461 39797 14473 39831
rect 14507 39828 14519 39831
rect 15654 39828 15660 39840
rect 14507 39800 15660 39828
rect 14507 39797 14519 39800
rect 14461 39791 14519 39797
rect 15654 39788 15660 39800
rect 15712 39788 15718 39840
rect 16390 39788 16396 39840
rect 16448 39788 16454 39840
rect 18414 39788 18420 39840
rect 18472 39828 18478 39840
rect 18877 39831 18935 39837
rect 18877 39828 18889 39831
rect 18472 39800 18889 39828
rect 18472 39788 18478 39800
rect 18877 39797 18889 39800
rect 18923 39797 18935 39831
rect 18877 39791 18935 39797
rect 1104 39738 28888 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 28888 39738
rect 1104 39664 28888 39686
rect 7006 39584 7012 39636
rect 7064 39584 7070 39636
rect 7653 39627 7711 39633
rect 7653 39593 7665 39627
rect 7699 39624 7711 39627
rect 8202 39624 8208 39636
rect 7699 39596 8208 39624
rect 7699 39593 7711 39596
rect 7653 39587 7711 39593
rect 8202 39584 8208 39596
rect 8260 39584 8266 39636
rect 9401 39627 9459 39633
rect 9401 39593 9413 39627
rect 9447 39624 9459 39627
rect 9674 39624 9680 39636
rect 9447 39596 9680 39624
rect 9447 39593 9459 39596
rect 9401 39587 9459 39593
rect 9674 39584 9680 39596
rect 9732 39584 9738 39636
rect 16025 39627 16083 39633
rect 16025 39593 16037 39627
rect 16071 39624 16083 39627
rect 16114 39624 16120 39636
rect 16071 39596 16120 39624
rect 16071 39593 16083 39596
rect 16025 39587 16083 39593
rect 16114 39584 16120 39596
rect 16172 39584 16178 39636
rect 10597 39559 10655 39565
rect 10597 39556 10609 39559
rect 8128 39528 10609 39556
rect 5534 39448 5540 39500
rect 5592 39488 5598 39500
rect 5629 39491 5687 39497
rect 5629 39488 5641 39491
rect 5592 39460 5641 39488
rect 5592 39448 5598 39460
rect 5629 39457 5641 39460
rect 5675 39457 5687 39491
rect 5629 39451 5687 39457
rect 7285 39491 7343 39497
rect 7285 39457 7297 39491
rect 7331 39488 7343 39491
rect 7650 39488 7656 39500
rect 7331 39460 7656 39488
rect 7331 39457 7343 39460
rect 7285 39451 7343 39457
rect 7650 39448 7656 39460
rect 7708 39448 7714 39500
rect 8128 39497 8156 39528
rect 10597 39525 10609 39528
rect 10643 39525 10655 39559
rect 10597 39519 10655 39525
rect 15013 39559 15071 39565
rect 15013 39525 15025 39559
rect 15059 39556 15071 39559
rect 15286 39556 15292 39568
rect 15059 39528 15292 39556
rect 15059 39525 15071 39528
rect 15013 39519 15071 39525
rect 15286 39516 15292 39528
rect 15344 39516 15350 39568
rect 8113 39491 8171 39497
rect 8113 39457 8125 39491
rect 8159 39457 8171 39491
rect 8113 39451 8171 39457
rect 9033 39491 9091 39497
rect 9033 39457 9045 39491
rect 9079 39488 9091 39491
rect 9677 39491 9735 39497
rect 9677 39488 9689 39491
rect 9079 39460 9689 39488
rect 9079 39457 9091 39460
rect 9033 39451 9091 39457
rect 9677 39457 9689 39460
rect 9723 39457 9735 39491
rect 9677 39451 9735 39457
rect 10870 39448 10876 39500
rect 10928 39488 10934 39500
rect 10928 39460 11008 39488
rect 10928 39448 10934 39460
rect 5902 39429 5908 39432
rect 5896 39420 5908 39429
rect 5863 39392 5908 39420
rect 5896 39383 5908 39392
rect 5902 39380 5908 39383
rect 5960 39380 5966 39432
rect 7469 39423 7527 39429
rect 7469 39420 7481 39423
rect 7300 39392 7481 39420
rect 7300 39364 7328 39392
rect 7469 39389 7481 39392
rect 7515 39389 7527 39423
rect 7469 39383 7527 39389
rect 9214 39380 9220 39432
rect 9272 39380 9278 39432
rect 10229 39423 10287 39429
rect 10229 39389 10241 39423
rect 10275 39389 10287 39423
rect 10229 39383 10287 39389
rect 7282 39312 7288 39364
rect 7340 39312 7346 39364
rect 7834 39312 7840 39364
rect 7892 39352 7898 39364
rect 10244 39352 10272 39383
rect 10778 39380 10784 39432
rect 10836 39380 10842 39432
rect 10980 39429 11008 39460
rect 11422 39448 11428 39500
rect 11480 39488 11486 39500
rect 11609 39491 11667 39497
rect 11609 39488 11621 39491
rect 11480 39460 11621 39488
rect 11480 39448 11486 39460
rect 11609 39457 11621 39460
rect 11655 39457 11667 39491
rect 11609 39451 11667 39457
rect 12066 39448 12072 39500
rect 12124 39448 12130 39500
rect 15105 39491 15163 39497
rect 15105 39457 15117 39491
rect 15151 39488 15163 39491
rect 18509 39491 18567 39497
rect 15151 39460 15424 39488
rect 15151 39457 15163 39460
rect 15105 39451 15163 39457
rect 10965 39423 11023 39429
rect 10965 39389 10977 39423
rect 11011 39389 11023 39423
rect 10965 39383 11023 39389
rect 11149 39423 11207 39429
rect 11149 39389 11161 39423
rect 11195 39389 11207 39423
rect 11149 39383 11207 39389
rect 11977 39423 12035 39429
rect 11977 39389 11989 39423
rect 12023 39420 12035 39423
rect 13630 39420 13636 39432
rect 12023 39392 13636 39420
rect 12023 39389 12035 39392
rect 11977 39383 12035 39389
rect 7892 39324 10272 39352
rect 7892 39312 7898 39324
rect 10686 39312 10692 39364
rect 10744 39352 10750 39364
rect 10873 39355 10931 39361
rect 10873 39352 10885 39355
rect 10744 39324 10885 39352
rect 10744 39312 10750 39324
rect 10873 39321 10885 39324
rect 10919 39321 10931 39355
rect 10873 39315 10931 39321
rect 8662 39244 8668 39296
rect 8720 39244 8726 39296
rect 9030 39244 9036 39296
rect 9088 39284 9094 39296
rect 11164 39284 11192 39383
rect 13630 39380 13636 39392
rect 13688 39380 13694 39432
rect 15396 39429 15424 39460
rect 18509 39457 18521 39491
rect 18555 39488 18567 39491
rect 19518 39488 19524 39500
rect 18555 39460 19524 39488
rect 18555 39457 18567 39460
rect 18509 39451 18567 39457
rect 19518 39448 19524 39460
rect 19576 39448 19582 39500
rect 15381 39423 15439 39429
rect 15381 39389 15393 39423
rect 15427 39389 15439 39423
rect 15381 39383 15439 39389
rect 15470 39380 15476 39432
rect 15528 39380 15534 39432
rect 15654 39380 15660 39432
rect 15712 39380 15718 39432
rect 15838 39380 15844 39432
rect 15896 39429 15902 39432
rect 15896 39420 15904 39429
rect 15896 39392 16344 39420
rect 15896 39383 15904 39392
rect 15896 39380 15902 39383
rect 14645 39355 14703 39361
rect 14645 39321 14657 39355
rect 14691 39352 14703 39355
rect 15194 39352 15200 39364
rect 14691 39324 15200 39352
rect 14691 39321 14703 39324
rect 14645 39315 14703 39321
rect 15194 39312 15200 39324
rect 15252 39352 15258 39364
rect 15562 39352 15568 39364
rect 15252 39324 15568 39352
rect 15252 39312 15258 39324
rect 15562 39312 15568 39324
rect 15620 39312 15626 39364
rect 15749 39355 15807 39361
rect 15749 39321 15761 39355
rect 15795 39352 15807 39355
rect 16022 39352 16028 39364
rect 15795 39324 16028 39352
rect 15795 39321 15807 39324
rect 15749 39315 15807 39321
rect 16022 39312 16028 39324
rect 16080 39312 16086 39364
rect 16316 39352 16344 39392
rect 16390 39380 16396 39432
rect 16448 39380 16454 39432
rect 18414 39420 18420 39432
rect 16500 39392 18420 39420
rect 16500 39364 16528 39392
rect 18414 39380 18420 39392
rect 18472 39380 18478 39432
rect 18690 39380 18696 39432
rect 18748 39380 18754 39432
rect 18877 39423 18935 39429
rect 18877 39389 18889 39423
rect 18923 39420 18935 39423
rect 19889 39423 19947 39429
rect 19889 39420 19901 39423
rect 18923 39392 19901 39420
rect 18923 39389 18935 39392
rect 18877 39383 18935 39389
rect 19889 39389 19901 39392
rect 19935 39389 19947 39423
rect 19889 39383 19947 39389
rect 16482 39352 16488 39364
rect 16316 39324 16488 39352
rect 16482 39312 16488 39324
rect 16540 39312 16546 39364
rect 9088 39256 11192 39284
rect 9088 39244 9094 39256
rect 16850 39244 16856 39296
rect 16908 39284 16914 39296
rect 17681 39287 17739 39293
rect 17681 39284 17693 39287
rect 16908 39256 17693 39284
rect 16908 39244 16914 39256
rect 17681 39253 17693 39256
rect 17727 39253 17739 39287
rect 17681 39247 17739 39253
rect 19150 39244 19156 39296
rect 19208 39284 19214 39296
rect 19337 39287 19395 39293
rect 19337 39284 19349 39287
rect 19208 39256 19349 39284
rect 19208 39244 19214 39256
rect 19337 39253 19349 39256
rect 19383 39253 19395 39287
rect 19337 39247 19395 39253
rect 1104 39194 28888 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 28888 39194
rect 1104 39120 28888 39142
rect 7742 39040 7748 39092
rect 7800 39040 7806 39092
rect 8113 39083 8171 39089
rect 8113 39049 8125 39083
rect 8159 39080 8171 39083
rect 10778 39080 10784 39092
rect 8159 39052 10784 39080
rect 8159 39049 8171 39052
rect 8113 39043 8171 39049
rect 10778 39040 10784 39052
rect 10836 39040 10842 39092
rect 13170 39040 13176 39092
rect 13228 39040 13234 39092
rect 17862 39040 17868 39092
rect 17920 39040 17926 39092
rect 18690 39040 18696 39092
rect 18748 39080 18754 39092
rect 20073 39083 20131 39089
rect 20073 39080 20085 39083
rect 18748 39052 20085 39080
rect 18748 39040 18754 39052
rect 20073 39049 20085 39052
rect 20119 39049 20131 39083
rect 20073 39043 20131 39049
rect 7561 39015 7619 39021
rect 7561 38981 7573 39015
rect 7607 39012 7619 39015
rect 8202 39012 8208 39024
rect 7607 38984 8208 39012
rect 7607 38981 7619 38984
rect 7561 38975 7619 38981
rect 8202 38972 8208 38984
rect 8260 38972 8266 39024
rect 8662 39021 8668 39024
rect 8656 39012 8668 39021
rect 8623 38984 8668 39012
rect 8656 38975 8668 38984
rect 8662 38972 8668 38975
rect 8720 38972 8726 39024
rect 19794 39012 19800 39024
rect 19720 38984 19800 39012
rect 7466 38904 7472 38956
rect 7524 38904 7530 38956
rect 7834 38904 7840 38956
rect 7892 38904 7898 38956
rect 8018 38904 8024 38956
rect 8076 38944 8082 38956
rect 8389 38947 8447 38953
rect 8389 38944 8401 38947
rect 8076 38916 8401 38944
rect 8076 38904 8082 38916
rect 8389 38913 8401 38916
rect 8435 38913 8447 38947
rect 9030 38944 9036 38956
rect 8389 38907 8447 38913
rect 8496 38916 9036 38944
rect 7929 38879 7987 38885
rect 7929 38845 7941 38879
rect 7975 38876 7987 38879
rect 8496 38876 8524 38916
rect 9030 38904 9036 38916
rect 9088 38904 9094 38956
rect 10502 38904 10508 38956
rect 10560 38944 10566 38956
rect 10965 38947 11023 38953
rect 10965 38944 10977 38947
rect 10560 38916 10977 38944
rect 10560 38904 10566 38916
rect 10965 38913 10977 38916
rect 11011 38913 11023 38947
rect 10965 38907 11023 38913
rect 11054 38904 11060 38956
rect 11112 38904 11118 38956
rect 12066 38904 12072 38956
rect 12124 38944 12130 38956
rect 12710 38944 12716 38956
rect 12124 38916 12716 38944
rect 12124 38904 12130 38916
rect 12710 38904 12716 38916
rect 12768 38944 12774 38956
rect 13357 38947 13415 38953
rect 13357 38944 13369 38947
rect 12768 38916 13369 38944
rect 12768 38904 12774 38916
rect 13357 38913 13369 38916
rect 13403 38913 13415 38947
rect 13357 38907 13415 38913
rect 13630 38904 13636 38956
rect 13688 38904 13694 38956
rect 13906 38904 13912 38956
rect 13964 38904 13970 38956
rect 14090 38904 14096 38956
rect 14148 38904 14154 38956
rect 15838 38904 15844 38956
rect 15896 38904 15902 38956
rect 15933 38947 15991 38953
rect 15933 38913 15945 38947
rect 15979 38913 15991 38947
rect 15933 38907 15991 38913
rect 16025 38947 16083 38953
rect 16025 38913 16037 38947
rect 16071 38944 16083 38947
rect 16298 38944 16304 38956
rect 16071 38916 16304 38944
rect 16071 38913 16083 38916
rect 16025 38907 16083 38913
rect 10594 38876 10600 38888
rect 7975 38848 8524 38876
rect 9784 38848 10600 38876
rect 7975 38845 7987 38848
rect 7929 38839 7987 38845
rect 9784 38817 9812 38848
rect 10594 38836 10600 38848
rect 10652 38836 10658 38888
rect 11072 38876 11100 38904
rect 11241 38879 11299 38885
rect 11241 38876 11253 38879
rect 11072 38848 11253 38876
rect 11241 38845 11253 38848
rect 11287 38876 11299 38879
rect 11882 38876 11888 38888
rect 11287 38848 11888 38876
rect 11287 38845 11299 38848
rect 11241 38839 11299 38845
rect 11882 38836 11888 38848
rect 11940 38836 11946 38888
rect 12802 38836 12808 38888
rect 12860 38836 12866 38888
rect 13170 38836 13176 38888
rect 13228 38876 13234 38888
rect 13648 38876 13676 38904
rect 14461 38879 14519 38885
rect 14461 38876 14473 38879
rect 13228 38848 14473 38876
rect 13228 38836 13234 38848
rect 14461 38845 14473 38848
rect 14507 38845 14519 38879
rect 14461 38839 14519 38845
rect 15105 38879 15163 38885
rect 15105 38845 15117 38879
rect 15151 38876 15163 38879
rect 15562 38876 15568 38888
rect 15151 38848 15568 38876
rect 15151 38845 15163 38848
rect 15105 38839 15163 38845
rect 15562 38836 15568 38848
rect 15620 38836 15626 38888
rect 15948 38876 15976 38907
rect 16298 38904 16304 38916
rect 16356 38904 16362 38956
rect 16850 38904 16856 38956
rect 16908 38904 16914 38956
rect 18989 38947 19047 38953
rect 18989 38913 19001 38947
rect 19035 38944 19047 38947
rect 19150 38944 19156 38956
rect 19035 38916 19156 38944
rect 19035 38913 19047 38916
rect 18989 38907 19047 38913
rect 19150 38904 19156 38916
rect 19208 38904 19214 38956
rect 19518 38904 19524 38956
rect 19576 38904 19582 38956
rect 19720 38953 19748 38984
rect 19794 38972 19800 38984
rect 19852 39012 19858 39024
rect 20441 39015 20499 39021
rect 20441 39012 20453 39015
rect 19852 38984 20453 39012
rect 19852 38972 19858 38984
rect 20441 38981 20453 38984
rect 20487 38981 20499 39015
rect 20441 38975 20499 38981
rect 19705 38947 19763 38953
rect 19705 38913 19717 38947
rect 19751 38913 19763 38947
rect 19705 38907 19763 38913
rect 19978 38904 19984 38956
rect 20036 38904 20042 38956
rect 20162 38904 20168 38956
rect 20220 38944 20226 38956
rect 20809 38947 20867 38953
rect 20809 38944 20821 38947
rect 20220 38916 20821 38944
rect 20220 38904 20226 38916
rect 20809 38913 20821 38916
rect 20855 38913 20867 38947
rect 20809 38907 20867 38913
rect 18138 38876 18144 38888
rect 15948 38848 18144 38876
rect 18138 38836 18144 38848
rect 18196 38836 18202 38888
rect 19245 38879 19303 38885
rect 19245 38845 19257 38879
rect 19291 38845 19303 38879
rect 19245 38839 19303 38845
rect 9769 38811 9827 38817
rect 9769 38777 9781 38811
rect 9815 38777 9827 38811
rect 9769 38771 9827 38777
rect 11057 38811 11115 38817
rect 11057 38777 11069 38811
rect 11103 38808 11115 38811
rect 12526 38808 12532 38820
rect 11103 38780 12532 38808
rect 11103 38777 11115 38780
rect 11057 38771 11115 38777
rect 12526 38768 12532 38780
rect 12584 38768 12590 38820
rect 13541 38811 13599 38817
rect 13541 38808 13553 38811
rect 13004 38780 13553 38808
rect 10042 38700 10048 38752
rect 10100 38700 10106 38752
rect 11149 38743 11207 38749
rect 11149 38709 11161 38743
rect 11195 38740 11207 38743
rect 11790 38740 11796 38752
rect 11195 38712 11796 38740
rect 11195 38709 11207 38712
rect 11149 38703 11207 38709
rect 11790 38700 11796 38712
rect 11848 38700 11854 38752
rect 12158 38700 12164 38752
rect 12216 38740 12222 38752
rect 12253 38743 12311 38749
rect 12253 38740 12265 38743
rect 12216 38712 12265 38740
rect 12216 38700 12222 38712
rect 12253 38709 12265 38712
rect 12299 38709 12311 38743
rect 12253 38703 12311 38709
rect 12342 38700 12348 38752
rect 12400 38740 12406 38752
rect 13004 38740 13032 38780
rect 13541 38777 13553 38780
rect 13587 38777 13599 38811
rect 13541 38771 13599 38777
rect 12400 38712 13032 38740
rect 12400 38700 12406 38712
rect 13998 38700 14004 38752
rect 14056 38700 14062 38752
rect 15378 38700 15384 38752
rect 15436 38740 15442 38752
rect 15657 38743 15715 38749
rect 15657 38740 15669 38743
rect 15436 38712 15669 38740
rect 15436 38700 15442 38712
rect 15657 38709 15669 38712
rect 15703 38709 15715 38743
rect 15657 38703 15715 38709
rect 17586 38700 17592 38752
rect 17644 38740 17650 38752
rect 18230 38740 18236 38752
rect 17644 38712 18236 38740
rect 17644 38700 17650 38712
rect 18230 38700 18236 38712
rect 18288 38740 18294 38752
rect 19260 38740 19288 38839
rect 18288 38712 19288 38740
rect 18288 38700 18294 38712
rect 19518 38700 19524 38752
rect 19576 38700 19582 38752
rect 20824 38740 20852 38907
rect 23106 38740 23112 38752
rect 20824 38712 23112 38740
rect 23106 38700 23112 38712
rect 23164 38700 23170 38752
rect 1104 38650 28888 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 28888 38650
rect 1104 38576 28888 38598
rect 9030 38496 9036 38548
rect 9088 38496 9094 38548
rect 9214 38496 9220 38548
rect 9272 38536 9278 38548
rect 9582 38536 9588 38548
rect 9272 38508 9588 38536
rect 9272 38496 9278 38508
rect 9582 38496 9588 38508
rect 9640 38536 9646 38548
rect 9677 38539 9735 38545
rect 9677 38536 9689 38539
rect 9640 38508 9689 38536
rect 9640 38496 9646 38508
rect 9677 38505 9689 38508
rect 9723 38505 9735 38539
rect 12710 38536 12716 38548
rect 9677 38499 9735 38505
rect 11440 38508 12716 38536
rect 11054 38428 11060 38480
rect 11112 38428 11118 38480
rect 9401 38403 9459 38409
rect 9401 38369 9413 38403
rect 9447 38400 9459 38403
rect 10042 38400 10048 38412
rect 9447 38372 10048 38400
rect 9447 38369 9459 38372
rect 9401 38363 9459 38369
rect 10042 38360 10048 38372
rect 10100 38360 10106 38412
rect 1210 38292 1216 38344
rect 1268 38332 1274 38344
rect 1489 38335 1547 38341
rect 1489 38332 1501 38335
rect 1268 38304 1501 38332
rect 1268 38292 1274 38304
rect 1489 38301 1501 38304
rect 1535 38332 1547 38335
rect 1949 38335 2007 38341
rect 1949 38332 1961 38335
rect 1535 38304 1961 38332
rect 1535 38301 1547 38304
rect 1489 38295 1547 38301
rect 1949 38301 1961 38304
rect 1995 38301 2007 38335
rect 1949 38295 2007 38301
rect 7282 38292 7288 38344
rect 7340 38332 7346 38344
rect 9217 38335 9275 38341
rect 9217 38332 9229 38335
rect 7340 38304 9229 38332
rect 7340 38292 7346 38304
rect 9217 38301 9229 38304
rect 9263 38332 9275 38335
rect 9263 38304 10456 38332
rect 9263 38301 9275 38304
rect 9217 38295 9275 38301
rect 1670 38156 1676 38208
rect 1728 38156 1734 38208
rect 10318 38156 10324 38208
rect 10376 38156 10382 38208
rect 10428 38196 10456 38304
rect 10502 38292 10508 38344
rect 10560 38292 10566 38344
rect 10781 38335 10839 38341
rect 10781 38301 10793 38335
rect 10827 38332 10839 38335
rect 11440 38332 11468 38508
rect 12710 38496 12716 38508
rect 12768 38496 12774 38548
rect 16850 38536 16856 38548
rect 14200 38508 16856 38536
rect 14200 38409 14228 38508
rect 16850 38496 16856 38508
rect 16908 38496 16914 38548
rect 17129 38539 17187 38545
rect 17129 38505 17141 38539
rect 17175 38505 17187 38539
rect 17129 38499 17187 38505
rect 17313 38539 17371 38545
rect 17313 38505 17325 38539
rect 17359 38536 17371 38539
rect 19334 38536 19340 38548
rect 17359 38508 19340 38536
rect 17359 38505 17371 38508
rect 17313 38499 17371 38505
rect 15562 38428 15568 38480
rect 15620 38428 15626 38480
rect 17144 38468 17172 38499
rect 19334 38496 19340 38508
rect 19392 38536 19398 38548
rect 19978 38536 19984 38548
rect 19392 38508 19984 38536
rect 19392 38496 19398 38508
rect 19978 38496 19984 38508
rect 20036 38496 20042 38548
rect 16776 38440 17172 38468
rect 18969 38471 19027 38477
rect 12437 38403 12495 38409
rect 12437 38369 12449 38403
rect 12483 38400 12495 38403
rect 14185 38403 14243 38409
rect 14185 38400 14197 38403
rect 12483 38372 14197 38400
rect 12483 38369 12495 38372
rect 12437 38363 12495 38369
rect 14185 38369 14197 38372
rect 14231 38369 14243 38403
rect 14185 38363 14243 38369
rect 15286 38360 15292 38412
rect 15344 38400 15350 38412
rect 16482 38400 16488 38412
rect 15344 38372 16488 38400
rect 15344 38360 15350 38372
rect 16482 38360 16488 38372
rect 16540 38400 16546 38412
rect 16776 38400 16804 38440
rect 18969 38437 18981 38471
rect 19015 38468 19027 38471
rect 19015 38440 19380 38468
rect 19015 38437 19027 38440
rect 18969 38431 19027 38437
rect 16540 38372 16804 38400
rect 16540 38360 16546 38372
rect 16850 38360 16856 38412
rect 16908 38400 16914 38412
rect 17586 38400 17592 38412
rect 16908 38372 17592 38400
rect 16908 38360 16914 38372
rect 17586 38360 17592 38372
rect 17644 38360 17650 38412
rect 19352 38409 19380 38440
rect 19337 38403 19395 38409
rect 19337 38369 19349 38403
rect 19383 38369 19395 38403
rect 19337 38363 19395 38369
rect 10827 38304 11468 38332
rect 10827 38301 10839 38304
rect 10781 38295 10839 38301
rect 12158 38292 12164 38344
rect 12216 38341 12222 38344
rect 12216 38332 12228 38341
rect 12805 38335 12863 38341
rect 12216 38304 12261 38332
rect 12216 38295 12228 38304
rect 12805 38301 12817 38335
rect 12851 38332 12863 38335
rect 12894 38332 12900 38344
rect 12851 38304 12900 38332
rect 12851 38301 12863 38304
rect 12805 38295 12863 38301
rect 12216 38292 12222 38295
rect 10689 38267 10747 38273
rect 10689 38233 10701 38267
rect 10735 38264 10747 38267
rect 12342 38264 12348 38276
rect 10735 38236 12348 38264
rect 10735 38233 10747 38236
rect 10689 38227 10747 38233
rect 12342 38224 12348 38236
rect 12400 38224 12406 38276
rect 12250 38196 12256 38208
rect 10428 38168 12256 38196
rect 12250 38156 12256 38168
rect 12308 38196 12314 38208
rect 12820 38196 12848 38295
rect 12894 38292 12900 38304
rect 12952 38292 12958 38344
rect 12989 38335 13047 38341
rect 12989 38301 13001 38335
rect 13035 38301 13047 38335
rect 12989 38295 13047 38301
rect 13004 38264 13032 38295
rect 13078 38292 13084 38344
rect 13136 38292 13142 38344
rect 13170 38292 13176 38344
rect 13228 38292 13234 38344
rect 13998 38332 14004 38344
rect 13280 38304 14004 38332
rect 13280 38264 13308 38304
rect 13998 38292 14004 38304
rect 14056 38292 14062 38344
rect 15838 38292 15844 38344
rect 15896 38292 15902 38344
rect 16025 38335 16083 38341
rect 16025 38301 16037 38335
rect 16071 38332 16083 38335
rect 16206 38332 16212 38344
rect 16071 38304 16212 38332
rect 16071 38301 16083 38304
rect 16025 38295 16083 38301
rect 16206 38292 16212 38304
rect 16264 38292 16270 38344
rect 16758 38332 16764 38344
rect 16500 38304 16764 38332
rect 13004 38236 13308 38264
rect 13449 38267 13507 38273
rect 13449 38233 13461 38267
rect 13495 38264 13507 38267
rect 14430 38267 14488 38273
rect 14430 38264 14442 38267
rect 13495 38236 14442 38264
rect 13495 38233 13507 38236
rect 13449 38227 13507 38233
rect 14430 38233 14442 38236
rect 14476 38233 14488 38267
rect 14430 38227 14488 38233
rect 16114 38224 16120 38276
rect 16172 38264 16178 38276
rect 16500 38273 16528 38304
rect 16758 38292 16764 38304
rect 16816 38332 16822 38344
rect 19794 38332 19800 38344
rect 16816 38304 19800 38332
rect 16816 38292 16822 38304
rect 19794 38292 19800 38304
rect 19852 38292 19858 38344
rect 16485 38267 16543 38273
rect 16485 38264 16497 38267
rect 16172 38236 16497 38264
rect 16172 38224 16178 38236
rect 16485 38233 16497 38236
rect 16531 38233 16543 38267
rect 16485 38227 16543 38233
rect 16574 38224 16580 38276
rect 16632 38264 16638 38276
rect 16945 38267 17003 38273
rect 16945 38264 16957 38267
rect 16632 38236 16957 38264
rect 16632 38224 16638 38236
rect 16945 38233 16957 38236
rect 16991 38233 17003 38267
rect 16945 38227 17003 38233
rect 17161 38267 17219 38273
rect 17161 38233 17173 38267
rect 17207 38264 17219 38267
rect 17856 38267 17914 38273
rect 17207 38236 17816 38264
rect 17207 38233 17219 38236
rect 17161 38227 17219 38233
rect 17788 38208 17816 38236
rect 17856 38233 17868 38267
rect 17902 38264 17914 38267
rect 18598 38264 18604 38276
rect 17902 38236 18604 38264
rect 17902 38233 17914 38236
rect 17856 38227 17914 38233
rect 18598 38224 18604 38236
rect 18656 38224 18662 38276
rect 12308 38168 12848 38196
rect 12308 38156 12314 38168
rect 15654 38156 15660 38208
rect 15712 38196 15718 38208
rect 15933 38199 15991 38205
rect 15933 38196 15945 38199
rect 15712 38168 15945 38196
rect 15712 38156 15718 38168
rect 15933 38165 15945 38168
rect 15979 38165 15991 38199
rect 15933 38159 15991 38165
rect 17770 38156 17776 38208
rect 17828 38156 17834 38208
rect 19886 38156 19892 38208
rect 19944 38196 19950 38208
rect 19981 38199 20039 38205
rect 19981 38196 19993 38199
rect 19944 38168 19993 38196
rect 19944 38156 19950 38168
rect 19981 38165 19993 38168
rect 20027 38165 20039 38199
rect 19981 38159 20039 38165
rect 1104 38106 28888 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 28888 38106
rect 1104 38032 28888 38054
rect 9030 37952 9036 38004
rect 9088 37952 9094 38004
rect 10502 37952 10508 38004
rect 10560 37992 10566 38004
rect 10873 37995 10931 38001
rect 10873 37992 10885 37995
rect 10560 37964 10885 37992
rect 10560 37952 10566 37964
rect 10873 37961 10885 37964
rect 10919 37961 10931 37995
rect 10873 37955 10931 37961
rect 12253 37995 12311 38001
rect 12253 37961 12265 37995
rect 12299 37992 12311 37995
rect 12802 37992 12808 38004
rect 12299 37964 12808 37992
rect 12299 37961 12311 37964
rect 12253 37955 12311 37961
rect 12802 37952 12808 37964
rect 12860 37952 12866 38004
rect 13078 37952 13084 38004
rect 13136 37992 13142 38004
rect 13449 37995 13507 38001
rect 13449 37992 13461 37995
rect 13136 37964 13461 37992
rect 13136 37952 13142 37964
rect 13449 37961 13461 37964
rect 13495 37992 13507 37995
rect 14090 37992 14096 38004
rect 13495 37964 14096 37992
rect 13495 37961 13507 37964
rect 13449 37955 13507 37961
rect 14090 37952 14096 37964
rect 14148 37952 14154 38004
rect 15013 37995 15071 38001
rect 15013 37992 15025 37995
rect 14384 37964 15025 37992
rect 5442 37924 5448 37936
rect 3160 37896 5448 37924
rect 1670 37816 1676 37868
rect 1728 37856 1734 37868
rect 3160 37865 3188 37896
rect 5442 37884 5448 37896
rect 5500 37924 5506 37936
rect 9048 37924 9076 37952
rect 9186 37927 9244 37933
rect 9186 37924 9198 37927
rect 5500 37896 6914 37924
rect 9048 37896 9198 37924
rect 5500 37884 5506 37896
rect 2685 37859 2743 37865
rect 2685 37856 2697 37859
rect 1728 37828 2697 37856
rect 1728 37816 1734 37828
rect 2685 37825 2697 37828
rect 2731 37825 2743 37859
rect 2685 37819 2743 37825
rect 3145 37859 3203 37865
rect 3145 37825 3157 37859
rect 3191 37825 3203 37859
rect 3401 37859 3459 37865
rect 3401 37856 3413 37859
rect 3145 37819 3203 37825
rect 3252 37828 3413 37856
rect 2501 37791 2559 37797
rect 2501 37757 2513 37791
rect 2547 37757 2559 37791
rect 2501 37751 2559 37757
rect 2869 37791 2927 37797
rect 2869 37757 2881 37791
rect 2915 37788 2927 37791
rect 3252 37788 3280 37828
rect 3401 37825 3413 37828
rect 3447 37825 3459 37859
rect 3401 37819 3459 37825
rect 2915 37760 3280 37788
rect 5077 37791 5135 37797
rect 2915 37757 2927 37760
rect 2869 37751 2927 37757
rect 5077 37757 5089 37791
rect 5123 37788 5135 37791
rect 5350 37788 5356 37800
rect 5123 37760 5356 37788
rect 5123 37757 5135 37760
rect 5077 37751 5135 37757
rect 2516 37652 2544 37751
rect 4525 37723 4583 37729
rect 4525 37689 4537 37723
rect 4571 37720 4583 37723
rect 5092 37720 5120 37751
rect 5350 37748 5356 37760
rect 5408 37748 5414 37800
rect 6886 37788 6914 37896
rect 9186 37893 9198 37896
rect 9232 37893 9244 37927
rect 9186 37887 9244 37893
rect 9582 37884 9588 37936
rect 9640 37924 9646 37936
rect 12986 37924 12992 37936
rect 9640 37896 12992 37924
rect 9640 37884 9646 37896
rect 8665 37859 8723 37865
rect 8665 37825 8677 37859
rect 8711 37856 8723 37859
rect 9030 37856 9036 37868
rect 8711 37828 9036 37856
rect 8711 37825 8723 37828
rect 8665 37819 8723 37825
rect 9030 37816 9036 37828
rect 9088 37816 9094 37868
rect 11057 37859 11115 37865
rect 11057 37825 11069 37859
rect 11103 37856 11115 37859
rect 11146 37856 11152 37868
rect 11103 37828 11152 37856
rect 11103 37825 11115 37828
rect 11057 37819 11115 37825
rect 11146 37816 11152 37828
rect 11204 37816 11210 37868
rect 11238 37816 11244 37868
rect 11296 37816 11302 37868
rect 11624 37865 11652 37896
rect 12986 37884 12992 37896
rect 13044 37924 13050 37936
rect 14384 37933 14412 37964
rect 15013 37961 15025 37964
rect 15059 37961 15071 37995
rect 15013 37955 15071 37961
rect 16393 37995 16451 38001
rect 16393 37961 16405 37995
rect 16439 37992 16451 37995
rect 16439 37964 18276 37992
rect 16439 37961 16451 37964
rect 16393 37955 16451 37961
rect 13725 37927 13783 37933
rect 13725 37924 13737 37927
rect 13044 37896 13737 37924
rect 13044 37884 13050 37896
rect 13725 37893 13737 37896
rect 13771 37893 13783 37927
rect 13725 37887 13783 37893
rect 14369 37927 14427 37933
rect 14369 37893 14381 37927
rect 14415 37893 14427 37927
rect 14369 37887 14427 37893
rect 14734 37884 14740 37936
rect 14792 37924 14798 37936
rect 15289 37927 15347 37933
rect 15289 37924 15301 37927
rect 14792 37896 15301 37924
rect 14792 37884 14798 37896
rect 15289 37893 15301 37896
rect 15335 37893 15347 37927
rect 15289 37887 15347 37893
rect 15378 37884 15384 37936
rect 15436 37884 15442 37936
rect 16114 37884 16120 37936
rect 16172 37884 16178 37936
rect 11609 37859 11667 37865
rect 11609 37825 11621 37859
rect 11655 37825 11667 37859
rect 11609 37819 11667 37825
rect 11790 37816 11796 37868
rect 11848 37816 11854 37868
rect 11882 37816 11888 37868
rect 11940 37816 11946 37868
rect 11977 37859 12035 37865
rect 11977 37825 11989 37859
rect 12023 37856 12035 37859
rect 12342 37856 12348 37868
rect 12023 37828 12348 37856
rect 12023 37825 12035 37828
rect 11977 37819 12035 37825
rect 12342 37816 12348 37828
rect 12400 37816 12406 37868
rect 14182 37816 14188 37868
rect 14240 37816 14246 37868
rect 14458 37816 14464 37868
rect 14516 37816 14522 37868
rect 15194 37865 15200 37868
rect 14553 37859 14611 37865
rect 14553 37825 14565 37859
rect 14599 37825 14611 37859
rect 15192 37856 15200 37865
rect 15155 37828 15200 37856
rect 14553 37819 14611 37825
rect 15192 37819 15200 37828
rect 7006 37788 7012 37800
rect 6886 37760 7012 37788
rect 7006 37748 7012 37760
rect 7064 37788 7070 37800
rect 8018 37788 8024 37800
rect 7064 37760 8024 37788
rect 7064 37748 7070 37760
rect 7282 37720 7288 37732
rect 4571 37692 5120 37720
rect 5184 37692 7288 37720
rect 4571 37689 4583 37692
rect 4525 37683 4583 37689
rect 4798 37652 4804 37664
rect 2516 37624 4804 37652
rect 4798 37612 4804 37624
rect 4856 37652 4862 37664
rect 5184 37652 5212 37692
rect 7282 37680 7288 37692
rect 7340 37680 7346 37732
rect 7392 37729 7420 37760
rect 8018 37748 8024 37760
rect 8076 37788 8082 37800
rect 8941 37791 8999 37797
rect 8941 37788 8953 37791
rect 8076 37760 8953 37788
rect 8076 37748 8082 37760
rect 8941 37757 8953 37760
rect 8987 37757 8999 37791
rect 11900 37788 11928 37816
rect 12618 37788 12624 37800
rect 11900 37760 12624 37788
rect 8941 37751 8999 37757
rect 12618 37748 12624 37760
rect 12676 37788 12682 37800
rect 12805 37791 12863 37797
rect 12805 37788 12817 37791
rect 12676 37760 12817 37788
rect 12676 37748 12682 37760
rect 12805 37757 12817 37760
rect 12851 37757 12863 37791
rect 14568 37788 14596 37819
rect 15194 37816 15200 37819
rect 15252 37816 15258 37868
rect 15562 37816 15568 37868
rect 15620 37816 15626 37868
rect 15654 37816 15660 37868
rect 15712 37816 15718 37868
rect 18248 37865 18276 37964
rect 18598 37952 18604 38004
rect 18656 37952 18662 38004
rect 19426 37952 19432 38004
rect 19484 37992 19490 38004
rect 19521 37995 19579 38001
rect 19521 37992 19533 37995
rect 19484 37964 19533 37992
rect 19484 37952 19490 37964
rect 19521 37961 19533 37964
rect 19567 37961 19579 37995
rect 19521 37955 19579 37961
rect 16393 37859 16451 37865
rect 16393 37825 16405 37859
rect 16439 37856 16451 37859
rect 18233 37859 18291 37865
rect 16439 37828 17908 37856
rect 16439 37825 16451 37828
rect 16393 37819 16451 37825
rect 17880 37800 17908 37828
rect 18233 37825 18245 37859
rect 18279 37825 18291 37859
rect 19705 37859 19763 37865
rect 19705 37856 19717 37859
rect 18233 37819 18291 37825
rect 18340 37828 19717 37856
rect 15930 37788 15936 37800
rect 14568 37760 15936 37788
rect 12805 37751 12863 37757
rect 15930 37748 15936 37760
rect 15988 37748 15994 37800
rect 17310 37748 17316 37800
rect 17368 37748 17374 37800
rect 17862 37748 17868 37800
rect 17920 37788 17926 37800
rect 18340 37788 18368 37828
rect 19705 37825 19717 37828
rect 19751 37825 19763 37859
rect 19705 37819 19763 37825
rect 17920 37760 18368 37788
rect 17920 37748 17926 37760
rect 18414 37748 18420 37800
rect 18472 37788 18478 37800
rect 19153 37791 19211 37797
rect 19153 37788 19165 37791
rect 18472 37760 19165 37788
rect 18472 37748 18478 37760
rect 19153 37757 19165 37760
rect 19199 37757 19211 37791
rect 19153 37751 19211 37757
rect 19886 37748 19892 37800
rect 19944 37748 19950 37800
rect 7377 37723 7435 37729
rect 7377 37689 7389 37723
rect 7423 37689 7435 37723
rect 7377 37683 7435 37689
rect 14737 37723 14795 37729
rect 14737 37689 14749 37723
rect 14783 37720 14795 37723
rect 15470 37720 15476 37732
rect 14783 37692 15476 37720
rect 14783 37689 14795 37692
rect 14737 37683 14795 37689
rect 15470 37680 15476 37692
rect 15528 37680 15534 37732
rect 16301 37723 16359 37729
rect 16301 37689 16313 37723
rect 16347 37720 16359 37723
rect 16761 37723 16819 37729
rect 16761 37720 16773 37723
rect 16347 37692 16773 37720
rect 16347 37689 16359 37692
rect 16301 37683 16359 37689
rect 16761 37689 16773 37692
rect 16807 37689 16819 37723
rect 16761 37683 16819 37689
rect 4856 37624 5212 37652
rect 4856 37612 4862 37624
rect 5626 37612 5632 37664
rect 5684 37612 5690 37664
rect 10321 37655 10379 37661
rect 10321 37621 10333 37655
rect 10367 37652 10379 37655
rect 10502 37652 10508 37664
rect 10367 37624 10508 37652
rect 10367 37621 10379 37624
rect 10321 37615 10379 37621
rect 10502 37612 10508 37624
rect 10560 37612 10566 37664
rect 17678 37612 17684 37664
rect 17736 37612 17742 37664
rect 1104 37562 28888 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 28888 37562
rect 1104 37488 28888 37510
rect 11146 37408 11152 37460
rect 11204 37448 11210 37460
rect 12434 37448 12440 37460
rect 11204 37420 12440 37448
rect 11204 37408 11210 37420
rect 12434 37408 12440 37420
rect 12492 37448 12498 37460
rect 12621 37451 12679 37457
rect 12621 37448 12633 37451
rect 12492 37420 12633 37448
rect 12492 37408 12498 37420
rect 12621 37417 12633 37420
rect 12667 37417 12679 37451
rect 12621 37411 12679 37417
rect 12894 37408 12900 37460
rect 12952 37448 12958 37460
rect 13725 37451 13783 37457
rect 13725 37448 13737 37451
rect 12952 37420 13737 37448
rect 12952 37408 12958 37420
rect 13725 37417 13737 37420
rect 13771 37417 13783 37451
rect 13725 37411 13783 37417
rect 14182 37408 14188 37460
rect 14240 37448 14246 37460
rect 14461 37451 14519 37457
rect 14461 37448 14473 37451
rect 14240 37420 14473 37448
rect 14240 37408 14246 37420
rect 14461 37417 14473 37420
rect 14507 37417 14519 37451
rect 14461 37411 14519 37417
rect 16482 37408 16488 37460
rect 16540 37448 16546 37460
rect 16540 37420 17724 37448
rect 16540 37408 16546 37420
rect 11422 37380 11428 37392
rect 10888 37352 11428 37380
rect 9030 37272 9036 37324
rect 9088 37272 9094 37324
rect 10888 37321 10916 37352
rect 11422 37340 11428 37352
rect 11480 37340 11486 37392
rect 13906 37380 13912 37392
rect 11716 37352 13912 37380
rect 10873 37315 10931 37321
rect 10873 37281 10885 37315
rect 10919 37281 10931 37315
rect 10873 37275 10931 37281
rect 11054 37272 11060 37324
rect 11112 37312 11118 37324
rect 11609 37315 11667 37321
rect 11609 37312 11621 37315
rect 11112 37284 11621 37312
rect 11112 37272 11118 37284
rect 11609 37281 11621 37284
rect 11655 37281 11667 37315
rect 11609 37275 11667 37281
rect 4985 37247 5043 37253
rect 4985 37213 4997 37247
rect 5031 37244 5043 37247
rect 5031 37216 5488 37244
rect 5031 37213 5043 37216
rect 4985 37207 5043 37213
rect 5460 37188 5488 37216
rect 7006 37204 7012 37256
rect 7064 37204 7070 37256
rect 10318 37204 10324 37256
rect 10376 37244 10382 37256
rect 10965 37247 11023 37253
rect 10965 37244 10977 37247
rect 10376 37216 10977 37244
rect 10376 37204 10382 37216
rect 10965 37213 10977 37216
rect 11011 37213 11023 37247
rect 10965 37207 11023 37213
rect 5258 37185 5264 37188
rect 5252 37139 5264 37185
rect 5258 37136 5264 37139
rect 5316 37136 5322 37188
rect 5442 37136 5448 37188
rect 5500 37136 5506 37188
rect 6362 37068 6368 37120
rect 6420 37068 6426 37120
rect 11333 37111 11391 37117
rect 11333 37077 11345 37111
rect 11379 37108 11391 37111
rect 11716 37108 11744 37352
rect 13906 37340 13912 37352
rect 13964 37340 13970 37392
rect 16209 37383 16267 37389
rect 16209 37349 16221 37383
rect 16255 37349 16267 37383
rect 16209 37343 16267 37349
rect 12253 37315 12311 37321
rect 12253 37281 12265 37315
rect 12299 37312 12311 37315
rect 12342 37312 12348 37324
rect 12299 37284 12348 37312
rect 12299 37281 12311 37284
rect 12253 37275 12311 37281
rect 12342 37272 12348 37284
rect 12400 37272 12406 37324
rect 12802 37272 12808 37324
rect 12860 37272 12866 37324
rect 14921 37315 14979 37321
rect 14921 37281 14933 37315
rect 14967 37312 14979 37315
rect 14967 37284 15424 37312
rect 14967 37281 14979 37284
rect 14921 37275 14979 37281
rect 12894 37204 12900 37256
rect 12952 37204 12958 37256
rect 13538 37204 13544 37256
rect 13596 37204 13602 37256
rect 14642 37204 14648 37256
rect 14700 37204 14706 37256
rect 14734 37204 14740 37256
rect 14792 37204 14798 37256
rect 15396 37253 15424 37284
rect 15013 37247 15071 37253
rect 15013 37213 15025 37247
rect 15059 37213 15071 37247
rect 15013 37207 15071 37213
rect 15381 37247 15439 37253
rect 15381 37213 15393 37247
rect 15427 37244 15439 37247
rect 16224 37244 16252 37343
rect 17586 37272 17592 37324
rect 17644 37272 17650 37324
rect 17696 37312 17724 37420
rect 17862 37408 17868 37460
rect 17920 37448 17926 37460
rect 18049 37451 18107 37457
rect 18049 37448 18061 37451
rect 17920 37420 18061 37448
rect 17920 37408 17926 37420
rect 18049 37417 18061 37420
rect 18095 37417 18107 37451
rect 18049 37411 18107 37417
rect 18414 37408 18420 37460
rect 18472 37408 18478 37460
rect 17957 37315 18015 37321
rect 17957 37312 17969 37315
rect 17696 37284 17969 37312
rect 17957 37281 17969 37284
rect 18003 37312 18015 37315
rect 19886 37312 19892 37324
rect 18003 37284 19892 37312
rect 18003 37281 18015 37284
rect 17957 37275 18015 37281
rect 19886 37272 19892 37284
rect 19944 37272 19950 37324
rect 15427 37216 16252 37244
rect 17333 37247 17391 37253
rect 15427 37213 15439 37216
rect 15381 37207 15439 37213
rect 17333 37213 17345 37247
rect 17379 37244 17391 37247
rect 17678 37244 17684 37256
rect 17379 37216 17684 37244
rect 17379 37213 17391 37216
rect 17333 37207 17391 37213
rect 12912 37176 12940 37204
rect 14458 37176 14464 37188
rect 12912 37148 14464 37176
rect 14458 37136 14464 37148
rect 14516 37176 14522 37188
rect 15028 37176 15056 37207
rect 17678 37204 17684 37216
rect 17736 37204 17742 37256
rect 18233 37247 18291 37253
rect 18233 37213 18245 37247
rect 18279 37244 18291 37247
rect 19518 37244 19524 37256
rect 18279 37216 19524 37244
rect 18279 37213 18291 37216
rect 18233 37207 18291 37213
rect 19518 37204 19524 37216
rect 19576 37204 19582 37256
rect 14516 37148 15056 37176
rect 14516 37136 14522 37148
rect 15930 37136 15936 37188
rect 15988 37136 15994 37188
rect 11379 37080 11744 37108
rect 11379 37077 11391 37080
rect 11333 37071 11391 37077
rect 1104 37018 28888 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 28888 37018
rect 1104 36944 28888 36966
rect 5077 36907 5135 36913
rect 5077 36873 5089 36907
rect 5123 36904 5135 36907
rect 5258 36904 5264 36916
rect 5123 36876 5264 36904
rect 5123 36873 5135 36876
rect 5077 36867 5135 36873
rect 5258 36864 5264 36876
rect 5316 36864 5322 36916
rect 12894 36864 12900 36916
rect 12952 36864 12958 36916
rect 14642 36864 14648 36916
rect 14700 36904 14706 36916
rect 15194 36904 15200 36916
rect 14700 36876 15200 36904
rect 14700 36864 14706 36876
rect 15194 36864 15200 36876
rect 15252 36904 15258 36916
rect 16574 36904 16580 36916
rect 15252 36876 16580 36904
rect 15252 36864 15258 36876
rect 12342 36796 12348 36848
rect 12400 36836 12406 36848
rect 12400 36808 13032 36836
rect 12400 36796 12406 36808
rect 4798 36728 4804 36780
rect 4856 36768 4862 36780
rect 5261 36771 5319 36777
rect 5261 36768 5273 36771
rect 4856 36740 5273 36768
rect 4856 36728 4862 36740
rect 5261 36737 5273 36740
rect 5307 36737 5319 36771
rect 5261 36731 5319 36737
rect 5445 36771 5503 36777
rect 5445 36737 5457 36771
rect 5491 36768 5503 36771
rect 5626 36768 5632 36780
rect 5491 36740 5632 36768
rect 5491 36737 5503 36740
rect 5445 36731 5503 36737
rect 5626 36728 5632 36740
rect 5684 36728 5690 36780
rect 11238 36728 11244 36780
rect 11296 36768 11302 36780
rect 11698 36768 11704 36780
rect 11296 36740 11704 36768
rect 11296 36728 11302 36740
rect 11698 36728 11704 36740
rect 11756 36768 11762 36780
rect 12253 36771 12311 36777
rect 12253 36768 12265 36771
rect 11756 36740 12265 36768
rect 11756 36728 11762 36740
rect 12253 36737 12265 36740
rect 12299 36737 12311 36771
rect 12253 36731 12311 36737
rect 12434 36728 12440 36780
rect 12492 36728 12498 36780
rect 13004 36777 13032 36808
rect 15672 36777 15700 36876
rect 16574 36864 16580 36876
rect 16632 36904 16638 36916
rect 16961 36907 17019 36913
rect 16961 36904 16973 36907
rect 16632 36876 16973 36904
rect 16632 36864 16638 36876
rect 16961 36873 16973 36876
rect 17007 36873 17019 36907
rect 16961 36867 17019 36873
rect 17129 36907 17187 36913
rect 17129 36873 17141 36907
rect 17175 36904 17187 36907
rect 17862 36904 17868 36916
rect 17175 36876 17868 36904
rect 17175 36873 17187 36876
rect 17129 36867 17187 36873
rect 17862 36864 17868 36876
rect 17920 36864 17926 36916
rect 15749 36839 15807 36845
rect 15749 36805 15761 36839
rect 15795 36836 15807 36839
rect 16206 36836 16212 36848
rect 15795 36808 16212 36836
rect 15795 36805 15807 36808
rect 15749 36799 15807 36805
rect 16206 36796 16212 36808
rect 16264 36836 16270 36848
rect 16761 36839 16819 36845
rect 16761 36836 16773 36839
rect 16264 36808 16773 36836
rect 16264 36796 16270 36808
rect 16761 36805 16773 36808
rect 16807 36805 16819 36839
rect 16761 36799 16819 36805
rect 12989 36771 13047 36777
rect 12989 36737 13001 36771
rect 13035 36737 13047 36771
rect 12989 36731 13047 36737
rect 15657 36771 15715 36777
rect 15657 36737 15669 36771
rect 15703 36737 15715 36771
rect 15657 36731 15715 36737
rect 15930 36728 15936 36780
rect 15988 36728 15994 36780
rect 6362 36660 6368 36712
rect 6420 36700 6426 36712
rect 7009 36703 7067 36709
rect 7009 36700 7021 36703
rect 6420 36672 7021 36700
rect 6420 36660 6426 36672
rect 7009 36669 7021 36672
rect 7055 36669 7067 36703
rect 7009 36663 7067 36669
rect 12437 36635 12495 36641
rect 12437 36601 12449 36635
rect 12483 36632 12495 36635
rect 12526 36632 12532 36644
rect 12483 36604 12532 36632
rect 12483 36601 12495 36604
rect 12437 36595 12495 36601
rect 12526 36592 12532 36604
rect 12584 36592 12590 36644
rect 15933 36635 15991 36641
rect 15933 36601 15945 36635
rect 15979 36632 15991 36635
rect 17310 36632 17316 36644
rect 15979 36604 17316 36632
rect 15979 36601 15991 36604
rect 15933 36595 15991 36601
rect 17310 36592 17316 36604
rect 17368 36592 17374 36644
rect 5626 36524 5632 36576
rect 5684 36564 5690 36576
rect 6457 36567 6515 36573
rect 6457 36564 6469 36567
rect 5684 36536 6469 36564
rect 5684 36524 5690 36536
rect 6457 36533 6469 36536
rect 6503 36533 6515 36567
rect 6457 36527 6515 36533
rect 16022 36524 16028 36576
rect 16080 36564 16086 36576
rect 16945 36567 17003 36573
rect 16945 36564 16957 36567
rect 16080 36536 16957 36564
rect 16080 36524 16086 36536
rect 16945 36533 16957 36536
rect 16991 36533 17003 36567
rect 16945 36527 17003 36533
rect 1104 36474 28888 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 28888 36474
rect 1104 36400 28888 36422
rect 5261 36159 5319 36165
rect 5261 36125 5273 36159
rect 5307 36156 5319 36159
rect 5350 36156 5356 36168
rect 5307 36128 5356 36156
rect 5307 36125 5319 36128
rect 5261 36119 5319 36125
rect 5350 36116 5356 36128
rect 5408 36116 5414 36168
rect 6454 36116 6460 36168
rect 6512 36156 6518 36168
rect 7469 36159 7527 36165
rect 7469 36156 7481 36159
rect 6512 36128 7481 36156
rect 6512 36116 6518 36128
rect 7469 36125 7481 36128
rect 7515 36125 7527 36159
rect 7469 36119 7527 36125
rect 5534 36097 5540 36100
rect 5528 36051 5540 36097
rect 5534 36048 5540 36051
rect 5592 36048 5598 36100
rect 4798 35980 4804 36032
rect 4856 36020 4862 36032
rect 4893 36023 4951 36029
rect 4893 36020 4905 36023
rect 4856 35992 4905 36020
rect 4856 35980 4862 35992
rect 4893 35989 4905 35992
rect 4939 35989 4951 36023
rect 4893 35983 4951 35989
rect 6086 35980 6092 36032
rect 6144 36020 6150 36032
rect 6641 36023 6699 36029
rect 6641 36020 6653 36023
rect 6144 35992 6653 36020
rect 6144 35980 6150 35992
rect 6641 35989 6653 35992
rect 6687 35989 6699 36023
rect 6641 35983 6699 35989
rect 6914 35980 6920 36032
rect 6972 35980 6978 36032
rect 1104 35930 28888 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 28888 35930
rect 1104 35856 28888 35878
rect 4525 35819 4583 35825
rect 4525 35785 4537 35819
rect 4571 35816 4583 35819
rect 5534 35816 5540 35828
rect 4571 35788 5540 35816
rect 4571 35785 4583 35788
rect 4525 35779 4583 35785
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 6454 35776 6460 35828
rect 6512 35776 6518 35828
rect 16206 35776 16212 35828
rect 16264 35776 16270 35828
rect 16758 35776 16764 35828
rect 16816 35776 16822 35828
rect 5626 35748 5632 35760
rect 4908 35720 5632 35748
rect 3881 35683 3939 35689
rect 3881 35649 3893 35683
rect 3927 35680 3939 35683
rect 4341 35683 4399 35689
rect 4341 35680 4353 35683
rect 3927 35652 4353 35680
rect 3927 35649 3939 35652
rect 3881 35643 3939 35649
rect 4341 35649 4353 35652
rect 4387 35680 4399 35683
rect 4798 35680 4804 35692
rect 4387 35652 4804 35680
rect 4387 35649 4399 35652
rect 4341 35643 4399 35649
rect 4798 35640 4804 35652
rect 4856 35640 4862 35692
rect 4908 35689 4936 35720
rect 5626 35708 5632 35720
rect 5684 35708 5690 35760
rect 6914 35748 6920 35760
rect 5736 35720 6920 35748
rect 4893 35683 4951 35689
rect 4893 35649 4905 35683
rect 4939 35649 4951 35683
rect 4893 35643 4951 35649
rect 4982 35640 4988 35692
rect 5040 35680 5046 35692
rect 5534 35680 5540 35692
rect 5040 35652 5540 35680
rect 5040 35640 5046 35652
rect 5534 35640 5540 35652
rect 5592 35640 5598 35692
rect 4157 35615 4215 35621
rect 4157 35581 4169 35615
rect 4203 35612 4215 35615
rect 5736 35612 5764 35720
rect 6914 35708 6920 35720
rect 6972 35708 6978 35760
rect 16025 35751 16083 35757
rect 16025 35717 16037 35751
rect 16071 35748 16083 35751
rect 16776 35748 16804 35776
rect 16071 35720 16804 35748
rect 16071 35717 16083 35720
rect 16025 35711 16083 35717
rect 7570 35683 7628 35689
rect 7570 35680 7582 35683
rect 6840 35652 7582 35680
rect 4203 35584 5764 35612
rect 4203 35581 4215 35584
rect 4157 35575 4215 35581
rect 6086 35572 6092 35624
rect 6144 35612 6150 35624
rect 6546 35612 6552 35624
rect 6144 35584 6552 35612
rect 6144 35572 6150 35584
rect 6546 35572 6552 35584
rect 6604 35572 6610 35624
rect 5169 35547 5227 35553
rect 5169 35513 5181 35547
rect 5215 35544 5227 35547
rect 6840 35544 6868 35652
rect 7570 35649 7582 35652
rect 7616 35649 7628 35683
rect 7570 35643 7628 35649
rect 7837 35683 7895 35689
rect 7837 35649 7849 35683
rect 7883 35680 7895 35683
rect 8018 35680 8024 35692
rect 7883 35652 8024 35680
rect 7883 35649 7895 35652
rect 7837 35643 7895 35649
rect 8018 35640 8024 35652
rect 8076 35640 8082 35692
rect 16298 35640 16304 35692
rect 16356 35640 16362 35692
rect 5215 35516 6914 35544
rect 5215 35513 5227 35516
rect 5169 35507 5227 35513
rect 6886 35488 6914 35516
rect 5258 35436 5264 35488
rect 5316 35476 5322 35488
rect 5445 35479 5503 35485
rect 5445 35476 5457 35479
rect 5316 35448 5457 35476
rect 5316 35436 5322 35448
rect 5445 35445 5457 35448
rect 5491 35445 5503 35479
rect 5445 35439 5503 35445
rect 5534 35436 5540 35488
rect 5592 35476 5598 35488
rect 6086 35476 6092 35488
rect 5592 35448 6092 35476
rect 5592 35436 5598 35448
rect 6086 35436 6092 35448
rect 6144 35436 6150 35488
rect 6886 35448 6920 35488
rect 6914 35436 6920 35448
rect 6972 35436 6978 35488
rect 15102 35436 15108 35488
rect 15160 35476 15166 35488
rect 16025 35479 16083 35485
rect 16025 35476 16037 35479
rect 15160 35448 16037 35476
rect 15160 35436 15166 35448
rect 16025 35445 16037 35448
rect 16071 35445 16083 35479
rect 16025 35439 16083 35445
rect 1104 35386 28888 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 28888 35386
rect 1104 35312 28888 35334
rect 5350 35232 5356 35284
rect 5408 35272 5414 35284
rect 5408 35244 6776 35272
rect 5408 35232 5414 35244
rect 6362 35204 6368 35216
rect 5092 35176 6368 35204
rect 5092 35077 5120 35176
rect 6362 35164 6368 35176
rect 6420 35164 6426 35216
rect 5261 35139 5319 35145
rect 5261 35105 5273 35139
rect 5307 35136 5319 35139
rect 5534 35136 5540 35148
rect 5307 35108 5540 35136
rect 5307 35105 5319 35108
rect 5261 35099 5319 35105
rect 5534 35096 5540 35108
rect 5592 35096 5598 35148
rect 6641 35139 6699 35145
rect 6641 35136 6653 35139
rect 5644 35108 6653 35136
rect 5644 35077 5672 35108
rect 6641 35105 6653 35108
rect 6687 35105 6699 35139
rect 6641 35099 6699 35105
rect 5077 35071 5135 35077
rect 5077 35037 5089 35071
rect 5123 35037 5135 35071
rect 5077 35031 5135 35037
rect 5629 35071 5687 35077
rect 5629 35037 5641 35071
rect 5675 35037 5687 35071
rect 5629 35031 5687 35037
rect 5997 35071 6055 35077
rect 5997 35037 6009 35071
rect 6043 35068 6055 35071
rect 6457 35071 6515 35077
rect 6457 35068 6469 35071
rect 6043 35040 6469 35068
rect 6043 35037 6055 35040
rect 5997 35031 6055 35037
rect 6457 35037 6469 35040
rect 6503 35037 6515 35071
rect 6457 35031 6515 35037
rect 5353 35003 5411 35009
rect 5353 34969 5365 35003
rect 5399 35000 5411 35003
rect 5399 34972 5764 35000
rect 5399 34969 5411 34972
rect 5353 34963 5411 34969
rect 4893 34935 4951 34941
rect 4893 34901 4905 34935
rect 4939 34932 4951 34935
rect 5442 34932 5448 34944
rect 4939 34904 5448 34932
rect 4939 34901 4951 34904
rect 4893 34895 4951 34901
rect 5442 34892 5448 34904
rect 5500 34892 5506 34944
rect 5736 34932 5764 34972
rect 5810 34960 5816 35012
rect 5868 34960 5874 35012
rect 5902 34960 5908 35012
rect 5960 34960 5966 35012
rect 6656 35000 6684 35099
rect 6748 35077 6776 35244
rect 11698 35232 11704 35284
rect 11756 35232 11762 35284
rect 16390 35232 16396 35284
rect 16448 35272 16454 35284
rect 16945 35275 17003 35281
rect 16945 35272 16957 35275
rect 16448 35244 16957 35272
rect 16448 35232 16454 35244
rect 16945 35241 16957 35244
rect 16991 35241 17003 35275
rect 16945 35235 17003 35241
rect 6822 35164 6828 35216
rect 6880 35204 6886 35216
rect 14829 35207 14887 35213
rect 6880 35164 6914 35204
rect 14829 35173 14841 35207
rect 14875 35204 14887 35207
rect 16758 35204 16764 35216
rect 14875 35176 16764 35204
rect 14875 35173 14887 35176
rect 14829 35167 14887 35173
rect 16758 35164 16764 35176
rect 16816 35204 16822 35216
rect 17586 35204 17592 35216
rect 16816 35176 17592 35204
rect 16816 35164 16822 35176
rect 17586 35164 17592 35176
rect 17644 35204 17650 35216
rect 18049 35207 18107 35213
rect 18049 35204 18061 35207
rect 17644 35176 18061 35204
rect 17644 35164 17650 35176
rect 18049 35173 18061 35176
rect 18095 35173 18107 35207
rect 18049 35167 18107 35173
rect 6886 35136 6914 35164
rect 9677 35139 9735 35145
rect 9677 35136 9689 35139
rect 6886 35108 9689 35136
rect 6733 35071 6791 35077
rect 6733 35037 6745 35071
rect 6779 35037 6791 35071
rect 6733 35031 6791 35037
rect 7006 35028 7012 35080
rect 7064 35068 7070 35080
rect 9232 35077 9260 35108
rect 9677 35105 9689 35108
rect 9723 35136 9735 35139
rect 12986 35136 12992 35148
rect 9723 35108 12992 35136
rect 9723 35105 9735 35108
rect 9677 35099 9735 35105
rect 12986 35096 12992 35108
rect 13044 35096 13050 35148
rect 7101 35071 7159 35077
rect 7101 35068 7113 35071
rect 7064 35040 7113 35068
rect 7064 35028 7070 35040
rect 7101 35037 7113 35040
rect 7147 35037 7159 35071
rect 7101 35031 7159 35037
rect 9217 35071 9275 35077
rect 9217 35037 9229 35071
rect 9263 35037 9275 35071
rect 9217 35031 9275 35037
rect 9398 35028 9404 35080
rect 9456 35028 9462 35080
rect 11882 35028 11888 35080
rect 11940 35028 11946 35080
rect 12066 35028 12072 35080
rect 12124 35068 12130 35080
rect 12161 35071 12219 35077
rect 12161 35068 12173 35071
rect 12124 35040 12173 35068
rect 12124 35028 12130 35040
rect 12161 35037 12173 35040
rect 12207 35037 12219 35071
rect 12161 35031 12219 35037
rect 16574 35028 16580 35080
rect 16632 35028 16638 35080
rect 9033 35003 9091 35009
rect 9033 35000 9045 35003
rect 6012 34972 6500 35000
rect 6656 34972 9045 35000
rect 6012 34932 6040 34972
rect 6472 34944 6500 34972
rect 9033 34969 9045 34972
rect 9079 35000 9091 35003
rect 9122 35000 9128 35012
rect 9079 34972 9128 35000
rect 9079 34969 9091 34972
rect 9033 34963 9091 34969
rect 9122 34960 9128 34972
rect 9180 34960 9186 35012
rect 5736 34904 6040 34932
rect 6178 34892 6184 34944
rect 6236 34892 6242 34944
rect 6454 34892 6460 34944
rect 6512 34892 6518 34944
rect 6546 34892 6552 34944
rect 6604 34932 6610 34944
rect 6825 34935 6883 34941
rect 6825 34932 6837 34935
rect 6604 34904 6837 34932
rect 6604 34892 6610 34904
rect 6825 34901 6837 34904
rect 6871 34901 6883 34935
rect 6825 34895 6883 34901
rect 6914 34892 6920 34944
rect 6972 34932 6978 34944
rect 7009 34935 7067 34941
rect 7009 34932 7021 34935
rect 6972 34904 7021 34932
rect 6972 34892 6978 34904
rect 7009 34901 7021 34904
rect 7055 34901 7067 34935
rect 7009 34895 7067 34901
rect 12069 34935 12127 34941
rect 12069 34901 12081 34935
rect 12115 34932 12127 34935
rect 12342 34932 12348 34944
rect 12115 34904 12348 34932
rect 12115 34901 12127 34904
rect 12069 34895 12127 34901
rect 12342 34892 12348 34904
rect 12400 34892 12406 34944
rect 14918 34892 14924 34944
rect 14976 34932 14982 34944
rect 16025 34935 16083 34941
rect 16025 34932 16037 34935
rect 14976 34904 16037 34932
rect 14976 34892 14982 34904
rect 16025 34901 16037 34904
rect 16071 34932 16083 34935
rect 16298 34932 16304 34944
rect 16071 34904 16304 34932
rect 16071 34901 16083 34904
rect 16025 34895 16083 34901
rect 16298 34892 16304 34904
rect 16356 34892 16362 34944
rect 1104 34842 28888 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 28888 34842
rect 1104 34768 28888 34790
rect 5718 34688 5724 34740
rect 5776 34728 5782 34740
rect 6822 34728 6828 34740
rect 5776 34700 6828 34728
rect 5776 34688 5782 34700
rect 6822 34688 6828 34700
rect 6880 34688 6886 34740
rect 7006 34688 7012 34740
rect 7064 34688 7070 34740
rect 10594 34728 10600 34740
rect 9876 34700 10600 34728
rect 6178 34620 6184 34672
rect 6236 34660 6242 34672
rect 6236 34632 7328 34660
rect 6236 34620 6242 34632
rect 5077 34595 5135 34601
rect 5077 34561 5089 34595
rect 5123 34561 5135 34595
rect 5077 34555 5135 34561
rect 5092 34524 5120 34555
rect 5258 34552 5264 34604
rect 5316 34552 5322 34604
rect 5626 34552 5632 34604
rect 5684 34592 5690 34604
rect 6641 34595 6699 34601
rect 6641 34592 6653 34595
rect 5684 34564 6653 34592
rect 5684 34552 5690 34564
rect 6641 34561 6653 34564
rect 6687 34561 6699 34595
rect 6641 34555 6699 34561
rect 6730 34552 6736 34604
rect 6788 34552 6794 34604
rect 6822 34552 6828 34604
rect 6880 34552 6886 34604
rect 7300 34601 7328 34632
rect 9876 34604 9904 34700
rect 10594 34688 10600 34700
rect 10652 34688 10658 34740
rect 12986 34688 12992 34740
rect 13044 34688 13050 34740
rect 14277 34731 14335 34737
rect 14277 34697 14289 34731
rect 14323 34728 14335 34731
rect 14734 34728 14740 34740
rect 14323 34700 14740 34728
rect 14323 34697 14335 34700
rect 14277 34691 14335 34697
rect 14734 34688 14740 34700
rect 14792 34688 14798 34740
rect 16206 34728 16212 34740
rect 14936 34700 16212 34728
rect 10502 34620 10508 34672
rect 10560 34620 10566 34672
rect 10870 34660 10876 34672
rect 10612 34632 10876 34660
rect 7285 34595 7343 34601
rect 7285 34561 7297 34595
rect 7331 34561 7343 34595
rect 7285 34555 7343 34561
rect 8849 34595 8907 34601
rect 8849 34561 8861 34595
rect 8895 34592 8907 34595
rect 8895 34564 9720 34592
rect 8895 34561 8907 34564
rect 8849 34555 8907 34561
rect 9692 34536 9720 34564
rect 9858 34552 9864 34604
rect 9916 34552 9922 34604
rect 10045 34595 10103 34601
rect 10045 34561 10057 34595
rect 10091 34592 10103 34595
rect 10134 34592 10140 34604
rect 10091 34564 10140 34592
rect 10091 34561 10103 34564
rect 10045 34555 10103 34561
rect 10134 34552 10140 34564
rect 10192 34592 10198 34604
rect 10520 34592 10548 34620
rect 10192 34564 10548 34592
rect 10192 34552 10198 34564
rect 5537 34527 5595 34533
rect 5537 34524 5549 34527
rect 5092 34496 5549 34524
rect 5537 34493 5549 34496
rect 5583 34524 5595 34527
rect 5718 34524 5724 34536
rect 5583 34496 5724 34524
rect 5583 34493 5595 34496
rect 5537 34487 5595 34493
rect 5718 34484 5724 34496
rect 5776 34484 5782 34536
rect 6454 34484 6460 34536
rect 6512 34484 6518 34536
rect 9398 34484 9404 34536
rect 9456 34484 9462 34536
rect 9674 34484 9680 34536
rect 9732 34524 9738 34536
rect 9769 34527 9827 34533
rect 9769 34524 9781 34527
rect 9732 34496 9781 34524
rect 9732 34484 9738 34496
rect 9769 34493 9781 34496
rect 9815 34493 9827 34527
rect 9769 34487 9827 34493
rect 9950 34484 9956 34536
rect 10008 34484 10014 34536
rect 10229 34527 10287 34533
rect 10229 34493 10241 34527
rect 10275 34524 10287 34527
rect 10612 34524 10640 34632
rect 10870 34620 10876 34632
rect 10928 34660 10934 34672
rect 12069 34663 12127 34669
rect 12069 34660 12081 34663
rect 10928 34632 12081 34660
rect 10928 34620 10934 34632
rect 12069 34629 12081 34632
rect 12115 34629 12127 34663
rect 12069 34623 12127 34629
rect 12621 34663 12679 34669
rect 12621 34629 12633 34663
rect 12667 34660 12679 34663
rect 12802 34660 12808 34672
rect 12667 34632 12808 34660
rect 12667 34629 12679 34632
rect 12621 34623 12679 34629
rect 12802 34620 12808 34632
rect 12860 34620 12866 34672
rect 14936 34660 14964 34700
rect 16206 34688 16212 34700
rect 16264 34688 16270 34740
rect 14844 34632 14964 34660
rect 10689 34595 10747 34601
rect 10689 34561 10701 34595
rect 10735 34592 10747 34595
rect 10778 34592 10784 34604
rect 10735 34564 10784 34592
rect 10735 34561 10747 34564
rect 10689 34555 10747 34561
rect 10778 34552 10784 34564
rect 10836 34552 10842 34604
rect 12250 34552 12256 34604
rect 12308 34552 12314 34604
rect 14182 34552 14188 34604
rect 14240 34552 14246 34604
rect 14642 34552 14648 34604
rect 14700 34592 14706 34604
rect 14844 34601 14872 34632
rect 15378 34620 15384 34672
rect 15436 34660 15442 34672
rect 16390 34660 16396 34672
rect 15436 34632 16396 34660
rect 15436 34620 15442 34632
rect 16390 34620 16396 34632
rect 16448 34660 16454 34672
rect 16761 34663 16819 34669
rect 16761 34660 16773 34663
rect 16448 34632 16773 34660
rect 16448 34620 16454 34632
rect 16761 34629 16773 34632
rect 16807 34629 16819 34663
rect 16761 34623 16819 34629
rect 14829 34595 14887 34601
rect 14829 34592 14841 34595
rect 14700 34564 14841 34592
rect 14700 34552 14706 34564
rect 14829 34561 14841 34564
rect 14875 34561 14887 34595
rect 14829 34555 14887 34561
rect 14918 34552 14924 34604
rect 14976 34552 14982 34604
rect 15102 34552 15108 34604
rect 15160 34552 15166 34604
rect 15562 34552 15568 34604
rect 15620 34552 15626 34604
rect 10275 34496 10640 34524
rect 10873 34527 10931 34533
rect 10275 34493 10287 34496
rect 10229 34487 10287 34493
rect 10873 34493 10885 34527
rect 10919 34524 10931 34527
rect 11238 34524 11244 34536
rect 10919 34496 11244 34524
rect 10919 34493 10931 34496
rect 10873 34487 10931 34493
rect 11238 34484 11244 34496
rect 11296 34484 11302 34536
rect 19426 34484 19432 34536
rect 19484 34484 19490 34536
rect 9030 34416 9036 34468
rect 9088 34456 9094 34468
rect 15378 34456 15384 34468
rect 9088 34428 15384 34456
rect 9088 34416 9094 34428
rect 15378 34416 15384 34428
rect 15436 34416 15442 34468
rect 4890 34348 4896 34400
rect 4948 34348 4954 34400
rect 7926 34348 7932 34400
rect 7984 34348 7990 34400
rect 15286 34348 15292 34400
rect 15344 34348 15350 34400
rect 17862 34348 17868 34400
rect 17920 34388 17926 34400
rect 18049 34391 18107 34397
rect 18049 34388 18061 34391
rect 17920 34360 18061 34388
rect 17920 34348 17926 34360
rect 18049 34357 18061 34360
rect 18095 34357 18107 34391
rect 18049 34351 18107 34357
rect 18782 34348 18788 34400
rect 18840 34348 18846 34400
rect 1104 34298 28888 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 28888 34298
rect 1104 34224 28888 34246
rect 5626 34144 5632 34196
rect 5684 34144 5690 34196
rect 5810 34144 5816 34196
rect 5868 34184 5874 34196
rect 6365 34187 6423 34193
rect 6365 34184 6377 34187
rect 5868 34156 6377 34184
rect 5868 34144 5874 34156
rect 6365 34153 6377 34156
rect 6411 34153 6423 34187
rect 6365 34147 6423 34153
rect 8665 34187 8723 34193
rect 8665 34153 8677 34187
rect 8711 34184 8723 34187
rect 9674 34184 9680 34196
rect 8711 34156 9680 34184
rect 8711 34153 8723 34156
rect 8665 34147 8723 34153
rect 9674 34144 9680 34156
rect 9732 34144 9738 34196
rect 9950 34144 9956 34196
rect 10008 34184 10014 34196
rect 10413 34187 10471 34193
rect 10413 34184 10425 34187
rect 10008 34156 10425 34184
rect 10008 34144 10014 34156
rect 10413 34153 10425 34156
rect 10459 34153 10471 34187
rect 10413 34147 10471 34153
rect 12342 34144 12348 34196
rect 12400 34184 12406 34196
rect 15838 34184 15844 34196
rect 12400 34156 15844 34184
rect 12400 34144 12406 34156
rect 10965 34119 11023 34125
rect 10965 34085 10977 34119
rect 11011 34116 11023 34119
rect 12618 34116 12624 34128
rect 11011 34088 12624 34116
rect 11011 34085 11023 34088
rect 10965 34079 11023 34085
rect 12618 34076 12624 34088
rect 12676 34076 12682 34128
rect 5460 34020 7236 34048
rect 4249 33983 4307 33989
rect 4249 33949 4261 33983
rect 4295 33980 4307 33983
rect 5460 33980 5488 34020
rect 7208 33992 7236 34020
rect 4295 33952 5488 33980
rect 4295 33949 4307 33952
rect 4249 33943 4307 33949
rect 6914 33940 6920 33992
rect 6972 33940 6978 33992
rect 7190 33940 7196 33992
rect 7248 33980 7254 33992
rect 7285 33983 7343 33989
rect 7285 33980 7297 33983
rect 7248 33952 7297 33980
rect 7248 33940 7254 33952
rect 7285 33949 7297 33952
rect 7331 33980 7343 33983
rect 9033 33983 9091 33989
rect 9033 33980 9045 33983
rect 7331 33952 9045 33980
rect 7331 33949 7343 33952
rect 7285 33943 7343 33949
rect 9033 33949 9045 33952
rect 9079 33949 9091 33983
rect 9033 33943 9091 33949
rect 9122 33940 9128 33992
rect 9180 33980 9186 33992
rect 9289 33983 9347 33989
rect 9289 33980 9301 33983
rect 9180 33952 9301 33980
rect 9180 33940 9186 33952
rect 9289 33949 9301 33952
rect 9335 33949 9347 33983
rect 9289 33943 9347 33949
rect 10686 33940 10692 33992
rect 10744 33940 10750 33992
rect 11238 33940 11244 33992
rect 11296 33940 11302 33992
rect 11514 33940 11520 33992
rect 11572 33940 11578 33992
rect 12526 33940 12532 33992
rect 12584 33940 12590 33992
rect 12636 33989 12664 34076
rect 13096 34048 13124 34156
rect 15838 34144 15844 34156
rect 15896 34144 15902 34196
rect 16301 34187 16359 34193
rect 16301 34153 16313 34187
rect 16347 34184 16359 34187
rect 16574 34184 16580 34196
rect 16347 34156 16580 34184
rect 16347 34153 16359 34156
rect 16301 34147 16359 34153
rect 16574 34144 16580 34156
rect 16632 34144 16638 34196
rect 17773 34187 17831 34193
rect 17773 34153 17785 34187
rect 17819 34184 17831 34187
rect 18782 34184 18788 34196
rect 17819 34156 18788 34184
rect 17819 34153 17831 34156
rect 17773 34147 17831 34153
rect 18782 34144 18788 34156
rect 18840 34144 18846 34196
rect 13173 34051 13231 34057
rect 13173 34048 13185 34051
rect 13096 34020 13185 34048
rect 13173 34017 13185 34020
rect 13219 34017 13231 34051
rect 13173 34011 13231 34017
rect 17586 34008 17592 34060
rect 17644 34048 17650 34060
rect 17865 34051 17923 34057
rect 17865 34048 17877 34051
rect 17644 34020 17877 34048
rect 17644 34008 17650 34020
rect 17865 34017 17877 34020
rect 17911 34017 17923 34051
rect 17865 34011 17923 34017
rect 12621 33983 12679 33989
rect 12621 33949 12633 33983
rect 12667 33949 12679 33983
rect 12621 33943 12679 33949
rect 4516 33915 4574 33921
rect 4516 33881 4528 33915
rect 4562 33912 4574 33915
rect 4890 33912 4896 33924
rect 4562 33884 4896 33912
rect 4562 33881 4574 33884
rect 4516 33875 4574 33881
rect 4890 33872 4896 33884
rect 4948 33872 4954 33924
rect 7552 33915 7610 33921
rect 7552 33881 7564 33915
rect 7598 33912 7610 33915
rect 7926 33912 7932 33924
rect 7598 33884 7932 33912
rect 7598 33881 7610 33884
rect 7552 33875 7610 33881
rect 7926 33872 7932 33884
rect 7984 33872 7990 33924
rect 12636 33912 12664 33943
rect 12710 33940 12716 33992
rect 12768 33940 12774 33992
rect 12897 33983 12955 33989
rect 12897 33949 12909 33983
rect 12943 33980 12955 33983
rect 12986 33980 12992 33992
rect 12943 33952 12992 33980
rect 12943 33949 12955 33952
rect 12897 33943 12955 33949
rect 12986 33940 12992 33952
rect 13044 33940 13050 33992
rect 14366 33940 14372 33992
rect 14424 33980 14430 33992
rect 14461 33983 14519 33989
rect 14461 33980 14473 33983
rect 14424 33952 14473 33980
rect 14424 33940 14430 33952
rect 14461 33949 14473 33952
rect 14507 33949 14519 33983
rect 14461 33943 14519 33949
rect 14642 33940 14648 33992
rect 14700 33940 14706 33992
rect 14921 33983 14979 33989
rect 14921 33949 14933 33983
rect 14967 33980 14979 33983
rect 15010 33980 15016 33992
rect 14967 33952 15016 33980
rect 14967 33949 14979 33952
rect 14921 33943 14979 33949
rect 15010 33940 15016 33952
rect 15068 33980 15074 33992
rect 16761 33983 16819 33989
rect 16761 33980 16773 33983
rect 15068 33952 16773 33980
rect 15068 33940 15074 33952
rect 16761 33949 16773 33952
rect 16807 33980 16819 33983
rect 17678 33980 17684 33992
rect 16807 33952 17684 33980
rect 16807 33949 16819 33952
rect 16761 33943 16819 33949
rect 17678 33940 17684 33952
rect 17736 33940 17742 33992
rect 17957 33983 18015 33989
rect 17957 33949 17969 33983
rect 18003 33980 18015 33983
rect 18785 33983 18843 33989
rect 18785 33980 18797 33983
rect 18003 33952 18797 33980
rect 18003 33949 18015 33952
rect 17957 33943 18015 33949
rect 18785 33949 18797 33952
rect 18831 33949 18843 33983
rect 18785 33943 18843 33949
rect 19150 33940 19156 33992
rect 19208 33980 19214 33992
rect 19337 33983 19395 33989
rect 19337 33980 19349 33983
rect 19208 33952 19349 33980
rect 19208 33940 19214 33952
rect 19337 33949 19349 33952
rect 19383 33949 19395 33983
rect 19337 33943 19395 33949
rect 22186 33940 22192 33992
rect 22244 33940 22250 33992
rect 25038 33940 25044 33992
rect 25096 33940 25102 33992
rect 12802 33912 12808 33924
rect 12636 33884 12808 33912
rect 12802 33872 12808 33884
rect 12860 33872 12866 33924
rect 15188 33915 15246 33921
rect 15188 33881 15200 33915
rect 15234 33912 15246 33915
rect 15286 33912 15292 33924
rect 15234 33884 15292 33912
rect 15234 33881 15246 33884
rect 15188 33875 15246 33881
rect 15286 33872 15292 33884
rect 15344 33872 15350 33924
rect 17494 33872 17500 33924
rect 17552 33872 17558 33924
rect 17589 33915 17647 33921
rect 17589 33881 17601 33915
rect 17635 33912 17647 33915
rect 17635 33884 19380 33912
rect 17635 33881 17647 33884
rect 17589 33875 17647 33881
rect 19352 33856 19380 33884
rect 12253 33847 12311 33853
rect 12253 33813 12265 33847
rect 12299 33844 12311 33847
rect 12434 33844 12440 33856
rect 12299 33816 12440 33844
rect 12299 33813 12311 33816
rect 12253 33807 12311 33813
rect 12434 33804 12440 33816
rect 12492 33804 12498 33856
rect 13814 33804 13820 33856
rect 13872 33804 13878 33856
rect 14550 33804 14556 33856
rect 14608 33804 14614 33856
rect 18046 33804 18052 33856
rect 18104 33844 18110 33856
rect 18233 33847 18291 33853
rect 18233 33844 18245 33847
rect 18104 33816 18245 33844
rect 18104 33804 18110 33816
rect 18233 33813 18245 33816
rect 18279 33813 18291 33847
rect 18233 33807 18291 33813
rect 19334 33804 19340 33856
rect 19392 33804 19398 33856
rect 19978 33804 19984 33856
rect 20036 33804 20042 33856
rect 21542 33804 21548 33856
rect 21600 33844 21606 33856
rect 21637 33847 21695 33853
rect 21637 33844 21649 33847
rect 21600 33816 21649 33844
rect 21600 33804 21606 33816
rect 21637 33813 21649 33816
rect 21683 33813 21695 33847
rect 21637 33807 21695 33813
rect 24486 33804 24492 33856
rect 24544 33804 24550 33856
rect 1104 33754 28888 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 28888 33754
rect 1104 33680 28888 33702
rect 9030 33640 9036 33652
rect 7116 33612 9036 33640
rect 7116 33581 7144 33612
rect 9030 33600 9036 33612
rect 9088 33640 9094 33652
rect 9125 33643 9183 33649
rect 9125 33640 9137 33643
rect 9088 33612 9137 33640
rect 9088 33600 9094 33612
rect 9125 33609 9137 33612
rect 9171 33609 9183 33643
rect 9125 33603 9183 33609
rect 9950 33600 9956 33652
rect 10008 33640 10014 33652
rect 10045 33643 10103 33649
rect 10045 33640 10057 33643
rect 10008 33612 10057 33640
rect 10008 33600 10014 33612
rect 10045 33609 10057 33612
rect 10091 33609 10103 33643
rect 10045 33603 10103 33609
rect 11241 33643 11299 33649
rect 11241 33609 11253 33643
rect 11287 33640 11299 33643
rect 11514 33640 11520 33652
rect 11287 33612 11520 33640
rect 11287 33609 11299 33612
rect 11241 33603 11299 33609
rect 11514 33600 11520 33612
rect 11572 33600 11578 33652
rect 15562 33600 15568 33652
rect 15620 33640 15626 33652
rect 16393 33643 16451 33649
rect 16393 33640 16405 33643
rect 15620 33612 16405 33640
rect 15620 33600 15626 33612
rect 16393 33609 16405 33612
rect 16439 33609 16451 33643
rect 16393 33603 16451 33609
rect 19150 33600 19156 33652
rect 19208 33600 19214 33652
rect 19426 33600 19432 33652
rect 19484 33640 19490 33652
rect 19521 33643 19579 33649
rect 19521 33640 19533 33643
rect 19484 33612 19533 33640
rect 19484 33600 19490 33612
rect 19521 33609 19533 33612
rect 19567 33609 19579 33643
rect 19521 33603 19579 33609
rect 7101 33575 7159 33581
rect 7101 33541 7113 33575
rect 7147 33541 7159 33575
rect 7101 33535 7159 33541
rect 10134 33532 10140 33584
rect 10192 33581 10198 33584
rect 10192 33575 10220 33581
rect 10208 33541 10220 33575
rect 10192 33535 10220 33541
rect 10192 33532 10198 33535
rect 11698 33532 11704 33584
rect 11756 33572 11762 33584
rect 11882 33572 11888 33584
rect 11756 33544 11888 33572
rect 11756 33532 11762 33544
rect 11882 33532 11888 33544
rect 11940 33532 11946 33584
rect 14550 33532 14556 33584
rect 14608 33572 14614 33584
rect 15258 33575 15316 33581
rect 15258 33572 15270 33575
rect 14608 33544 15270 33572
rect 14608 33532 14614 33544
rect 15258 33541 15270 33544
rect 15304 33541 15316 33575
rect 17862 33572 17868 33584
rect 15258 33535 15316 33541
rect 17788 33544 17868 33572
rect 5626 33464 5632 33516
rect 5684 33504 5690 33516
rect 5997 33507 6055 33513
rect 5997 33504 6009 33507
rect 5684 33476 6009 33504
rect 5684 33464 5690 33476
rect 5997 33473 6009 33476
rect 6043 33473 6055 33507
rect 5997 33467 6055 33473
rect 9674 33464 9680 33516
rect 9732 33464 9738 33516
rect 9858 33464 9864 33516
rect 9916 33504 9922 33516
rect 9953 33507 10011 33513
rect 9953 33504 9965 33507
rect 9916 33476 9965 33504
rect 9916 33464 9922 33476
rect 9953 33473 9965 33476
rect 9999 33473 10011 33507
rect 9953 33467 10011 33473
rect 12434 33464 12440 33516
rect 12492 33464 12498 33516
rect 14001 33507 14059 33513
rect 14001 33473 14013 33507
rect 14047 33504 14059 33507
rect 14182 33504 14188 33516
rect 14047 33476 14188 33504
rect 14047 33473 14059 33476
rect 14001 33467 14059 33473
rect 14182 33464 14188 33476
rect 14240 33464 14246 33516
rect 14458 33464 14464 33516
rect 14516 33464 14522 33516
rect 15010 33464 15016 33516
rect 15068 33464 15074 33516
rect 17586 33464 17592 33516
rect 17644 33504 17650 33516
rect 17788 33513 17816 33544
rect 17862 33532 17868 33544
rect 17920 33572 17926 33584
rect 24388 33575 24446 33581
rect 17920 33544 24164 33572
rect 17920 33532 17926 33544
rect 18046 33513 18052 33516
rect 17773 33507 17831 33513
rect 17773 33504 17785 33507
rect 17644 33476 17785 33504
rect 17644 33464 17650 33476
rect 17773 33473 17785 33476
rect 17819 33473 17831 33507
rect 18040 33504 18052 33513
rect 18007 33476 18052 33504
rect 17773 33467 17831 33473
rect 18040 33467 18052 33476
rect 18046 33464 18052 33467
rect 18104 33464 18110 33516
rect 19429 33507 19487 33513
rect 19429 33473 19441 33507
rect 19475 33473 19487 33507
rect 19429 33467 19487 33473
rect 19613 33507 19671 33513
rect 19613 33473 19625 33507
rect 19659 33504 19671 33507
rect 19978 33504 19984 33516
rect 19659 33476 19984 33504
rect 19659 33473 19671 33476
rect 19613 33467 19671 33473
rect 10594 33396 10600 33448
rect 10652 33396 10658 33448
rect 13814 33396 13820 33448
rect 13872 33436 13878 33448
rect 14274 33436 14280 33448
rect 13872 33408 14280 33436
rect 13872 33396 13878 33408
rect 14274 33396 14280 33408
rect 14332 33436 14338 33448
rect 14737 33439 14795 33445
rect 14737 33436 14749 33439
rect 14332 33408 14749 33436
rect 14332 33396 14338 33408
rect 14737 33405 14749 33408
rect 14783 33405 14795 33439
rect 19444 33436 19472 33467
rect 19978 33464 19984 33476
rect 20036 33464 20042 33516
rect 21085 33507 21143 33513
rect 21085 33473 21097 33507
rect 21131 33504 21143 33507
rect 21361 33507 21419 33513
rect 21361 33504 21373 33507
rect 21131 33476 21373 33504
rect 21131 33473 21143 33476
rect 21085 33467 21143 33473
rect 21361 33473 21373 33476
rect 21407 33473 21419 33507
rect 21361 33467 21419 33473
rect 19702 33436 19708 33448
rect 19444 33408 19708 33436
rect 14737 33399 14795 33405
rect 19702 33396 19708 33408
rect 19760 33396 19766 33448
rect 12066 33328 12072 33380
rect 12124 33328 12130 33380
rect 12526 33328 12532 33380
rect 12584 33368 12590 33380
rect 13357 33371 13415 33377
rect 13357 33368 13369 33371
rect 12584 33340 13369 33368
rect 12584 33328 12590 33340
rect 13357 33337 13369 33340
rect 13403 33337 13415 33371
rect 13357 33331 13415 33337
rect 14090 33328 14096 33380
rect 14148 33368 14154 33380
rect 14645 33371 14703 33377
rect 14645 33368 14657 33371
rect 14148 33340 14657 33368
rect 14148 33328 14154 33340
rect 14645 33337 14657 33340
rect 14691 33337 14703 33371
rect 14645 33331 14703 33337
rect 5445 33303 5503 33309
rect 5445 33269 5457 33303
rect 5491 33300 5503 33303
rect 5534 33300 5540 33312
rect 5491 33272 5540 33300
rect 5491 33269 5503 33272
rect 5445 33263 5503 33269
rect 5534 33260 5540 33272
rect 5592 33260 5598 33312
rect 7190 33260 7196 33312
rect 7248 33300 7254 33312
rect 8389 33303 8447 33309
rect 8389 33300 8401 33303
rect 7248 33272 8401 33300
rect 7248 33260 7254 33272
rect 8389 33269 8401 33272
rect 8435 33269 8447 33303
rect 8389 33263 8447 33269
rect 10321 33303 10379 33309
rect 10321 33269 10333 33303
rect 10367 33300 10379 33303
rect 11054 33300 11060 33312
rect 10367 33272 11060 33300
rect 10367 33269 10379 33272
rect 10321 33263 10379 33269
rect 11054 33260 11060 33272
rect 11112 33260 11118 33312
rect 11882 33260 11888 33312
rect 11940 33300 11946 33312
rect 12161 33303 12219 33309
rect 12161 33300 12173 33303
rect 11940 33272 12173 33300
rect 11940 33260 11946 33272
rect 12161 33269 12173 33272
rect 12207 33269 12219 33303
rect 12161 33263 12219 33269
rect 13078 33260 13084 33312
rect 13136 33260 13142 33312
rect 13906 33260 13912 33312
rect 13964 33300 13970 33312
rect 14277 33303 14335 33309
rect 14277 33300 14289 33303
rect 13964 33272 14289 33300
rect 13964 33260 13970 33272
rect 14277 33269 14289 33272
rect 14323 33269 14335 33303
rect 21376 33300 21404 33467
rect 21542 33464 21548 33516
rect 21600 33464 21606 33516
rect 21928 33513 21956 33544
rect 21913 33507 21971 33513
rect 21913 33473 21925 33507
rect 21959 33473 21971 33507
rect 22169 33507 22227 33513
rect 22169 33504 22181 33507
rect 21913 33467 21971 33473
rect 22020 33476 22181 33504
rect 21453 33439 21511 33445
rect 21453 33405 21465 33439
rect 21499 33436 21511 33439
rect 22020 33436 22048 33476
rect 22169 33473 22181 33476
rect 22215 33473 22227 33507
rect 22169 33467 22227 33473
rect 23750 33464 23756 33516
rect 23808 33464 23814 33516
rect 24136 33445 24164 33544
rect 24388 33541 24400 33575
rect 24434 33572 24446 33575
rect 24486 33572 24492 33584
rect 24434 33544 24492 33572
rect 24434 33541 24446 33544
rect 24388 33535 24446 33541
rect 24486 33532 24492 33544
rect 24544 33532 24550 33584
rect 21499 33408 22048 33436
rect 24121 33439 24179 33445
rect 21499 33405 21511 33408
rect 21453 33399 21511 33405
rect 24121 33405 24133 33439
rect 24167 33405 24179 33439
rect 26329 33439 26387 33445
rect 26329 33436 26341 33439
rect 24121 33399 24179 33405
rect 26206 33408 26341 33436
rect 23566 33368 23572 33380
rect 22848 33340 23572 33368
rect 22848 33300 22876 33340
rect 23566 33328 23572 33340
rect 23624 33328 23630 33380
rect 21376 33272 22876 33300
rect 14277 33263 14335 33269
rect 23290 33260 23296 33312
rect 23348 33260 23354 33312
rect 23658 33260 23664 33312
rect 23716 33260 23722 33312
rect 24136 33300 24164 33399
rect 25501 33371 25559 33377
rect 25501 33337 25513 33371
rect 25547 33368 25559 33371
rect 26206 33368 26234 33408
rect 26329 33405 26341 33408
rect 26375 33405 26387 33439
rect 26329 33399 26387 33405
rect 25547 33340 26234 33368
rect 25547 33337 25559 33340
rect 25501 33331 25559 33337
rect 25314 33300 25320 33312
rect 24136 33272 25320 33300
rect 25314 33260 25320 33272
rect 25372 33260 25378 33312
rect 25682 33260 25688 33312
rect 25740 33300 25746 33312
rect 25777 33303 25835 33309
rect 25777 33300 25789 33303
rect 25740 33272 25789 33300
rect 25740 33260 25746 33272
rect 25777 33269 25789 33272
rect 25823 33269 25835 33303
rect 25777 33263 25835 33269
rect 1104 33210 28888 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 28888 33210
rect 1104 33136 28888 33158
rect 5721 33099 5779 33105
rect 5721 33065 5733 33099
rect 5767 33065 5779 33099
rect 5721 33059 5779 33065
rect 5905 33099 5963 33105
rect 5905 33065 5917 33099
rect 5951 33096 5963 33099
rect 6914 33096 6920 33108
rect 5951 33068 6920 33096
rect 5951 33065 5963 33068
rect 5905 33059 5963 33065
rect 5736 33028 5764 33059
rect 6914 33056 6920 33068
rect 6972 33056 6978 33108
rect 10778 33056 10784 33108
rect 10836 33096 10842 33108
rect 10873 33099 10931 33105
rect 10873 33096 10885 33099
rect 10836 33068 10885 33096
rect 10836 33056 10842 33068
rect 10873 33065 10885 33068
rect 10919 33065 10931 33099
rect 10873 33059 10931 33065
rect 12342 33056 12348 33108
rect 12400 33096 12406 33108
rect 12437 33099 12495 33105
rect 12437 33096 12449 33099
rect 12400 33068 12449 33096
rect 12400 33056 12406 33068
rect 12437 33065 12449 33068
rect 12483 33065 12495 33099
rect 12437 33059 12495 33065
rect 14458 33056 14464 33108
rect 14516 33056 14522 33108
rect 16301 33099 16359 33105
rect 16301 33065 16313 33099
rect 16347 33096 16359 33099
rect 16758 33096 16764 33108
rect 16347 33068 16764 33096
rect 16347 33065 16359 33068
rect 16301 33059 16359 33065
rect 16758 33056 16764 33068
rect 16816 33056 16822 33108
rect 17494 33056 17500 33108
rect 17552 33056 17558 33108
rect 19334 33056 19340 33108
rect 19392 33096 19398 33108
rect 19429 33099 19487 33105
rect 19429 33096 19441 33099
rect 19392 33068 19441 33096
rect 19392 33056 19398 33068
rect 19429 33065 19441 33068
rect 19475 33065 19487 33099
rect 19429 33059 19487 33065
rect 21729 33099 21787 33105
rect 21729 33065 21741 33099
rect 21775 33096 21787 33099
rect 22186 33096 22192 33108
rect 21775 33068 22192 33096
rect 21775 33065 21787 33068
rect 21729 33059 21787 33065
rect 22186 33056 22192 33068
rect 22244 33056 22250 33108
rect 23750 33056 23756 33108
rect 23808 33056 23814 33108
rect 6181 33031 6239 33037
rect 6181 33028 6193 33031
rect 5736 33000 6193 33028
rect 6181 32997 6193 33000
rect 6227 33028 6239 33031
rect 6730 33028 6736 33040
rect 6227 33000 6736 33028
rect 6227 32997 6239 33000
rect 6181 32991 6239 32997
rect 6730 32988 6736 33000
rect 6788 32988 6794 33040
rect 9585 33031 9643 33037
rect 9585 32997 9597 33031
rect 9631 33028 9643 33031
rect 10686 33028 10692 33040
rect 9631 33000 10692 33028
rect 9631 32997 9643 33000
rect 9585 32991 9643 32997
rect 10686 32988 10692 33000
rect 10744 32988 10750 33040
rect 15933 33031 15991 33037
rect 15933 32997 15945 33031
rect 15979 33028 15991 33031
rect 16482 33028 16488 33040
rect 15979 33000 16488 33028
rect 15979 32997 15991 33000
rect 15933 32991 15991 32997
rect 16482 32988 16488 33000
rect 16540 32988 16546 33040
rect 17865 33031 17923 33037
rect 17865 32997 17877 33031
rect 17911 33028 17923 33031
rect 18233 33031 18291 33037
rect 18233 33028 18245 33031
rect 17911 33000 18245 33028
rect 17911 32997 17923 33000
rect 17865 32991 17923 32997
rect 18233 32997 18245 33000
rect 18279 33028 18291 33031
rect 18279 33000 19564 33028
rect 18279 32997 18291 33000
rect 18233 32991 18291 32997
rect 5537 32963 5595 32969
rect 5537 32929 5549 32963
rect 5583 32960 5595 32963
rect 6822 32960 6828 32972
rect 5583 32932 6828 32960
rect 5583 32929 5595 32932
rect 5537 32923 5595 32929
rect 6822 32920 6828 32932
rect 6880 32920 6886 32972
rect 9309 32963 9367 32969
rect 9309 32929 9321 32963
rect 9355 32960 9367 32963
rect 9858 32960 9864 32972
rect 9355 32932 9864 32960
rect 9355 32929 9367 32932
rect 9309 32923 9367 32929
rect 9858 32920 9864 32932
rect 9916 32920 9922 32972
rect 9950 32920 9956 32972
rect 10008 32960 10014 32972
rect 10229 32963 10287 32969
rect 10229 32960 10241 32963
rect 10008 32932 10241 32960
rect 10008 32920 10014 32932
rect 10229 32929 10241 32932
rect 10275 32929 10287 32963
rect 10229 32923 10287 32929
rect 11882 32920 11888 32972
rect 11940 32920 11946 32972
rect 13814 32920 13820 32972
rect 13872 32960 13878 32972
rect 15010 32960 15016 32972
rect 13872 32932 15016 32960
rect 13872 32920 13878 32932
rect 15010 32920 15016 32932
rect 15068 32920 15074 32972
rect 18693 32963 18751 32969
rect 18693 32929 18705 32963
rect 18739 32960 18751 32963
rect 18874 32960 18880 32972
rect 18739 32932 18880 32960
rect 18739 32929 18751 32932
rect 18693 32923 18751 32929
rect 18874 32920 18880 32932
rect 18932 32920 18938 32972
rect 19260 32932 19472 32960
rect 5442 32852 5448 32904
rect 5500 32852 5506 32904
rect 5626 32852 5632 32904
rect 5684 32892 5690 32904
rect 5721 32895 5779 32901
rect 5721 32892 5733 32895
rect 5684 32864 5733 32892
rect 5684 32852 5690 32864
rect 5721 32861 5733 32864
rect 5767 32861 5779 32895
rect 5721 32855 5779 32861
rect 6454 32852 6460 32904
rect 6512 32892 6518 32904
rect 6733 32895 6791 32901
rect 6733 32892 6745 32895
rect 6512 32864 6745 32892
rect 6512 32852 6518 32864
rect 6733 32861 6745 32864
rect 6779 32861 6791 32895
rect 6733 32855 6791 32861
rect 9217 32895 9275 32901
rect 9217 32861 9229 32895
rect 9263 32892 9275 32895
rect 9398 32892 9404 32904
rect 9263 32864 9404 32892
rect 9263 32861 9275 32864
rect 9217 32855 9275 32861
rect 9398 32852 9404 32864
rect 9456 32852 9462 32904
rect 11793 32895 11851 32901
rect 11793 32861 11805 32895
rect 11839 32892 11851 32895
rect 12342 32892 12348 32904
rect 11839 32864 12348 32892
rect 11839 32861 11851 32864
rect 11793 32855 11851 32861
rect 12342 32852 12348 32864
rect 12400 32852 12406 32904
rect 13561 32895 13619 32901
rect 13561 32861 13573 32895
rect 13607 32892 13619 32895
rect 13906 32892 13912 32904
rect 13607 32864 13912 32892
rect 13607 32861 13619 32864
rect 13561 32855 13619 32861
rect 13906 32852 13912 32864
rect 13964 32852 13970 32904
rect 14090 32852 14096 32904
rect 14148 32892 14154 32904
rect 14185 32895 14243 32901
rect 14185 32892 14197 32895
rect 14148 32864 14197 32892
rect 14148 32852 14154 32864
rect 14185 32861 14197 32864
rect 14231 32861 14243 32895
rect 14185 32855 14243 32861
rect 14274 32852 14280 32904
rect 14332 32852 14338 32904
rect 15657 32895 15715 32901
rect 15657 32861 15669 32895
rect 15703 32892 15715 32895
rect 17678 32892 17684 32904
rect 15703 32864 17684 32892
rect 15703 32861 15715 32864
rect 15657 32855 15715 32861
rect 17678 32852 17684 32864
rect 17736 32852 17742 32904
rect 17957 32895 18015 32901
rect 17957 32861 17969 32895
rect 18003 32861 18015 32895
rect 17957 32855 18015 32861
rect 18601 32895 18659 32901
rect 18601 32861 18613 32895
rect 18647 32892 18659 32895
rect 19260 32892 19288 32932
rect 18647 32864 19288 32892
rect 19337 32895 19395 32901
rect 18647 32861 18659 32864
rect 18601 32855 18659 32861
rect 19337 32861 19349 32895
rect 19383 32861 19395 32895
rect 19337 32855 19395 32861
rect 7101 32827 7159 32833
rect 7101 32793 7113 32827
rect 7147 32824 7159 32827
rect 7190 32824 7196 32836
rect 7147 32796 7196 32824
rect 7147 32793 7159 32796
rect 7101 32787 7159 32793
rect 7190 32784 7196 32796
rect 7248 32784 7254 32836
rect 14366 32784 14372 32836
rect 14424 32824 14430 32836
rect 14461 32827 14519 32833
rect 14461 32824 14473 32827
rect 14424 32796 14473 32824
rect 14424 32784 14430 32796
rect 14461 32793 14473 32796
rect 14507 32824 14519 32827
rect 14829 32827 14887 32833
rect 14829 32824 14841 32827
rect 14507 32796 14841 32824
rect 14507 32793 14519 32796
rect 14461 32787 14519 32793
rect 14829 32793 14841 32796
rect 14875 32824 14887 32827
rect 15933 32827 15991 32833
rect 15933 32824 15945 32827
rect 14875 32796 15945 32824
rect 14875 32793 14887 32796
rect 14829 32787 14887 32793
rect 15933 32793 15945 32796
rect 15979 32824 15991 32827
rect 16758 32824 16764 32836
rect 15979 32796 16764 32824
rect 15979 32793 15991 32796
rect 15933 32787 15991 32793
rect 16758 32784 16764 32796
rect 16816 32824 16822 32836
rect 17770 32824 17776 32836
rect 16816 32796 17776 32824
rect 16816 32784 16822 32796
rect 17770 32784 17776 32796
rect 17828 32784 17834 32836
rect 17972 32824 18000 32855
rect 19352 32824 19380 32855
rect 17972 32796 19380 32824
rect 19444 32824 19472 32932
rect 19536 32901 19564 33000
rect 19702 32988 19708 33040
rect 19760 33028 19766 33040
rect 23842 33028 23848 33040
rect 19760 33000 23848 33028
rect 19760 32988 19766 33000
rect 21174 32920 21180 32972
rect 21232 32920 21238 32972
rect 22296 32969 22324 33000
rect 23842 32988 23848 33000
rect 23900 32988 23906 33040
rect 21453 32963 21511 32969
rect 21453 32929 21465 32963
rect 21499 32960 21511 32963
rect 22189 32963 22247 32969
rect 22189 32960 22201 32963
rect 21499 32932 22201 32960
rect 21499 32929 21511 32932
rect 21453 32923 21511 32929
rect 22189 32929 22201 32932
rect 22235 32929 22247 32963
rect 22189 32923 22247 32929
rect 22281 32963 22339 32969
rect 22281 32929 22293 32963
rect 22327 32929 22339 32963
rect 22281 32923 22339 32929
rect 23201 32963 23259 32969
rect 23201 32929 23213 32963
rect 23247 32960 23259 32963
rect 23290 32960 23296 32972
rect 23247 32932 23296 32960
rect 23247 32929 23259 32932
rect 23201 32923 23259 32929
rect 23290 32920 23296 32932
rect 23348 32920 23354 32972
rect 23382 32920 23388 32972
rect 23440 32960 23446 32972
rect 25685 32963 25743 32969
rect 25685 32960 25697 32963
rect 23440 32932 25697 32960
rect 23440 32920 23446 32932
rect 25685 32929 25697 32932
rect 25731 32929 25743 32963
rect 25685 32923 25743 32929
rect 19521 32895 19579 32901
rect 19521 32861 19533 32895
rect 19567 32892 19579 32895
rect 19702 32892 19708 32904
rect 19567 32864 19708 32892
rect 19567 32861 19579 32864
rect 19521 32855 19579 32861
rect 19702 32852 19708 32864
rect 19760 32852 19766 32904
rect 19978 32852 19984 32904
rect 20036 32852 20042 32904
rect 21085 32895 21143 32901
rect 21085 32861 21097 32895
rect 21131 32892 21143 32895
rect 21910 32892 21916 32904
rect 21131 32864 21916 32892
rect 21131 32861 21143 32864
rect 21085 32855 21143 32861
rect 21910 32852 21916 32864
rect 21968 32852 21974 32904
rect 22097 32895 22155 32901
rect 22097 32861 22109 32895
rect 22143 32892 22155 32895
rect 22370 32892 22376 32904
rect 22143 32864 22376 32892
rect 22143 32861 22155 32864
rect 22097 32855 22155 32861
rect 22370 32852 22376 32864
rect 22428 32892 22434 32904
rect 23658 32892 23664 32904
rect 22428 32864 23664 32892
rect 22428 32852 22434 32864
rect 23658 32852 23664 32864
rect 23716 32852 23722 32904
rect 25130 32852 25136 32904
rect 25188 32852 25194 32904
rect 25774 32852 25780 32904
rect 25832 32852 25838 32904
rect 19444 32796 19932 32824
rect 18616 32768 18644 32796
rect 12158 32716 12164 32768
rect 12216 32716 12222 32768
rect 15746 32716 15752 32768
rect 15804 32716 15810 32768
rect 18598 32716 18604 32768
rect 18656 32716 18662 32768
rect 19904 32765 19932 32796
rect 19889 32759 19947 32765
rect 19889 32725 19901 32759
rect 19935 32756 19947 32759
rect 20162 32756 20168 32768
rect 19935 32728 20168 32756
rect 19935 32725 19947 32728
rect 19889 32719 19947 32725
rect 20162 32716 20168 32728
rect 20220 32716 20226 32768
rect 23658 32716 23664 32768
rect 23716 32756 23722 32768
rect 24489 32759 24547 32765
rect 24489 32756 24501 32759
rect 23716 32728 24501 32756
rect 23716 32716 23722 32728
rect 24489 32725 24501 32728
rect 24535 32725 24547 32759
rect 24489 32719 24547 32725
rect 24670 32716 24676 32768
rect 24728 32756 24734 32768
rect 25409 32759 25467 32765
rect 25409 32756 25421 32759
rect 24728 32728 25421 32756
rect 24728 32716 24734 32728
rect 25409 32725 25421 32728
rect 25455 32725 25467 32759
rect 25409 32719 25467 32725
rect 1104 32666 28888 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 28888 32666
rect 1104 32592 28888 32614
rect 6454 32512 6460 32564
rect 6512 32512 6518 32564
rect 10045 32555 10103 32561
rect 10045 32521 10057 32555
rect 10091 32552 10103 32555
rect 10594 32552 10600 32564
rect 10091 32524 10600 32552
rect 10091 32521 10103 32524
rect 10045 32515 10103 32521
rect 10594 32512 10600 32524
rect 10652 32512 10658 32564
rect 11241 32555 11299 32561
rect 11241 32521 11253 32555
rect 11287 32552 11299 32555
rect 11698 32552 11704 32564
rect 11287 32524 11704 32552
rect 11287 32521 11299 32524
rect 11241 32515 11299 32521
rect 11698 32512 11704 32524
rect 11756 32512 11762 32564
rect 11977 32555 12035 32561
rect 11977 32521 11989 32555
rect 12023 32552 12035 32555
rect 12066 32552 12072 32564
rect 12023 32524 12072 32552
rect 12023 32521 12035 32524
rect 11977 32515 12035 32521
rect 12066 32512 12072 32524
rect 12124 32512 12130 32564
rect 12526 32552 12532 32564
rect 12176 32524 12532 32552
rect 5261 32487 5319 32493
rect 5261 32453 5273 32487
rect 5307 32484 5319 32487
rect 10134 32484 10140 32496
rect 5307 32456 5672 32484
rect 5307 32453 5319 32456
rect 5261 32447 5319 32453
rect 5534 32376 5540 32428
rect 5592 32376 5598 32428
rect 5644 32416 5672 32456
rect 9876 32456 10140 32484
rect 5718 32416 5724 32428
rect 5776 32425 5782 32428
rect 5776 32419 5799 32425
rect 5644 32388 5724 32416
rect 5718 32376 5724 32388
rect 5787 32416 5799 32419
rect 6638 32416 6644 32428
rect 5787 32388 6644 32416
rect 5787 32385 5799 32388
rect 5776 32379 5799 32385
rect 5776 32376 5782 32379
rect 6638 32376 6644 32388
rect 6696 32376 6702 32428
rect 7581 32419 7639 32425
rect 7581 32385 7593 32419
rect 7627 32416 7639 32419
rect 7926 32416 7932 32428
rect 7627 32388 7932 32416
rect 7627 32385 7639 32388
rect 7581 32379 7639 32385
rect 7926 32376 7932 32388
rect 7984 32376 7990 32428
rect 9876 32425 9904 32456
rect 10134 32444 10140 32456
rect 10192 32444 10198 32496
rect 10778 32444 10784 32496
rect 10836 32444 10842 32496
rect 10888 32456 11652 32484
rect 9861 32419 9919 32425
rect 9861 32385 9873 32419
rect 9907 32385 9919 32419
rect 9861 32379 9919 32385
rect 10045 32419 10103 32425
rect 10045 32385 10057 32419
rect 10091 32416 10103 32419
rect 10796 32416 10824 32444
rect 10888 32428 10916 32456
rect 10091 32388 10824 32416
rect 10091 32385 10103 32388
rect 10045 32379 10103 32385
rect 10870 32376 10876 32428
rect 10928 32376 10934 32428
rect 11624 32425 11652 32456
rect 11057 32419 11115 32425
rect 11057 32385 11069 32419
rect 11103 32385 11115 32419
rect 11057 32379 11115 32385
rect 11609 32419 11667 32425
rect 11609 32385 11621 32419
rect 11655 32385 11667 32419
rect 11609 32379 11667 32385
rect 11793 32419 11851 32425
rect 11793 32385 11805 32419
rect 11839 32416 11851 32419
rect 12176 32416 12204 32524
rect 12526 32512 12532 32524
rect 12584 32512 12590 32564
rect 15746 32512 15752 32564
rect 15804 32552 15810 32564
rect 16390 32552 16396 32564
rect 15804 32524 16396 32552
rect 15804 32512 15810 32524
rect 16390 32512 16396 32524
rect 16448 32552 16454 32564
rect 17405 32555 17463 32561
rect 17405 32552 17417 32555
rect 16448 32524 17417 32552
rect 16448 32512 16454 32524
rect 17405 32521 17417 32524
rect 17451 32521 17463 32555
rect 17405 32515 17463 32521
rect 17678 32512 17684 32564
rect 17736 32552 17742 32564
rect 19610 32552 19616 32564
rect 17736 32524 19616 32552
rect 17736 32512 17742 32524
rect 19610 32512 19616 32524
rect 19668 32512 19674 32564
rect 21910 32512 21916 32564
rect 21968 32512 21974 32564
rect 23842 32512 23848 32564
rect 23900 32512 23906 32564
rect 24213 32555 24271 32561
rect 24213 32521 24225 32555
rect 24259 32521 24271 32555
rect 24213 32515 24271 32521
rect 13814 32484 13820 32496
rect 12452 32456 13820 32484
rect 12452 32425 12480 32456
rect 13814 32444 13820 32456
rect 13872 32444 13878 32496
rect 17034 32444 17040 32496
rect 17092 32484 17098 32496
rect 17696 32484 17724 32512
rect 23382 32484 23388 32496
rect 17092 32456 17724 32484
rect 22940 32456 23388 32484
rect 17092 32444 17098 32456
rect 11839 32388 12204 32416
rect 12437 32419 12495 32425
rect 11839 32385 11851 32388
rect 11793 32379 11851 32385
rect 12437 32385 12449 32419
rect 12483 32385 12495 32419
rect 12437 32379 12495 32385
rect 12704 32419 12762 32425
rect 12704 32385 12716 32419
rect 12750 32416 12762 32419
rect 13078 32416 13084 32428
rect 12750 32388 13084 32416
rect 12750 32385 12762 32388
rect 12704 32379 12762 32385
rect 7837 32351 7895 32357
rect 7837 32317 7849 32351
rect 7883 32317 7895 32351
rect 7837 32311 7895 32317
rect 10781 32351 10839 32357
rect 10781 32317 10793 32351
rect 10827 32317 10839 32351
rect 11072 32348 11100 32379
rect 11808 32348 11836 32379
rect 13078 32376 13084 32388
rect 13136 32376 13142 32428
rect 15010 32376 15016 32428
rect 15068 32376 15074 32428
rect 15286 32425 15292 32428
rect 15280 32379 15292 32425
rect 15286 32376 15292 32379
rect 15344 32376 15350 32428
rect 18874 32376 18880 32428
rect 18932 32376 18938 32428
rect 19153 32419 19211 32425
rect 19153 32385 19165 32419
rect 19199 32416 19211 32419
rect 19978 32416 19984 32428
rect 19199 32388 19984 32416
rect 19199 32385 19211 32388
rect 19153 32379 19211 32385
rect 19978 32376 19984 32388
rect 20036 32376 20042 32428
rect 22281 32419 22339 32425
rect 22281 32385 22293 32419
rect 22327 32416 22339 32419
rect 22370 32416 22376 32428
rect 22327 32388 22376 32416
rect 22327 32385 22339 32388
rect 22281 32379 22339 32385
rect 22370 32376 22376 32388
rect 22428 32376 22434 32428
rect 22940 32425 22968 32456
rect 23382 32444 23388 32456
rect 23440 32444 23446 32496
rect 23937 32487 23995 32493
rect 23937 32453 23949 32487
rect 23983 32484 23995 32487
rect 24228 32484 24256 32515
rect 25130 32512 25136 32564
rect 25188 32512 25194 32564
rect 23983 32456 24256 32484
rect 23983 32453 23995 32456
rect 23937 32447 23995 32453
rect 22925 32419 22983 32425
rect 22925 32385 22937 32419
rect 22971 32385 22983 32419
rect 22925 32379 22983 32385
rect 23201 32419 23259 32425
rect 23201 32385 23213 32419
rect 23247 32416 23259 32419
rect 23290 32416 23296 32428
rect 23247 32388 23296 32416
rect 23247 32385 23259 32388
rect 23201 32379 23259 32385
rect 11072 32320 11836 32348
rect 16761 32351 16819 32357
rect 10781 32311 10839 32317
rect 16761 32317 16773 32351
rect 16807 32317 16819 32351
rect 16761 32311 16819 32317
rect 842 32172 848 32224
rect 900 32212 906 32224
rect 1489 32215 1547 32221
rect 1489 32212 1501 32215
rect 900 32184 1501 32212
rect 900 32172 906 32184
rect 1489 32181 1501 32184
rect 1535 32181 1547 32215
rect 1489 32175 1547 32181
rect 5626 32172 5632 32224
rect 5684 32212 5690 32224
rect 5905 32215 5963 32221
rect 5905 32212 5917 32215
rect 5684 32184 5917 32212
rect 5684 32172 5690 32184
rect 5905 32181 5917 32184
rect 5951 32181 5963 32215
rect 5905 32175 5963 32181
rect 7190 32172 7196 32224
rect 7248 32212 7254 32224
rect 7852 32212 7880 32311
rect 10796 32280 10824 32311
rect 11054 32280 11060 32292
rect 10796 32252 11060 32280
rect 11054 32240 11060 32252
rect 11112 32280 11118 32292
rect 13817 32283 13875 32289
rect 11112 32252 11836 32280
rect 11112 32240 11118 32252
rect 11808 32221 11836 32252
rect 13817 32249 13829 32283
rect 13863 32280 13875 32283
rect 14182 32280 14188 32292
rect 13863 32252 14188 32280
rect 13863 32249 13875 32252
rect 13817 32243 13875 32249
rect 14182 32240 14188 32252
rect 14240 32240 14246 32292
rect 16393 32283 16451 32289
rect 16393 32249 16405 32283
rect 16439 32280 16451 32283
rect 16776 32280 16804 32311
rect 21910 32308 21916 32360
rect 21968 32348 21974 32360
rect 22189 32351 22247 32357
rect 22189 32348 22201 32351
rect 21968 32320 22201 32348
rect 21968 32308 21974 32320
rect 22189 32317 22201 32320
rect 22235 32348 22247 32351
rect 22940 32348 22968 32379
rect 23290 32376 23296 32388
rect 23348 32376 23354 32428
rect 23658 32376 23664 32428
rect 23716 32376 23722 32428
rect 24210 32376 24216 32428
rect 24268 32416 24274 32428
rect 24581 32419 24639 32425
rect 24581 32416 24593 32419
rect 24268 32388 24593 32416
rect 24268 32376 24274 32388
rect 24581 32385 24593 32388
rect 24627 32385 24639 32419
rect 24581 32379 24639 32385
rect 25041 32419 25099 32425
rect 25041 32385 25053 32419
rect 25087 32385 25099 32419
rect 25041 32379 25099 32385
rect 25225 32419 25283 32425
rect 25225 32385 25237 32419
rect 25271 32416 25283 32419
rect 25682 32416 25688 32428
rect 25271 32388 25688 32416
rect 25271 32385 25283 32388
rect 25225 32379 25283 32385
rect 22235 32320 22968 32348
rect 22235 32317 22247 32320
rect 22189 32311 22247 32317
rect 23566 32308 23572 32360
rect 23624 32308 23630 32360
rect 24670 32308 24676 32360
rect 24728 32308 24734 32360
rect 16439 32252 16804 32280
rect 18693 32283 18751 32289
rect 16439 32249 16451 32252
rect 16393 32243 16451 32249
rect 18693 32249 18705 32283
rect 18739 32280 18751 32283
rect 19426 32280 19432 32292
rect 18739 32252 19432 32280
rect 18739 32249 18751 32252
rect 18693 32243 18751 32249
rect 19426 32240 19432 32252
rect 19484 32240 19490 32292
rect 23842 32240 23848 32292
rect 23900 32280 23906 32292
rect 25056 32280 25084 32379
rect 25682 32376 25688 32388
rect 25740 32376 25746 32428
rect 27062 32376 27068 32428
rect 27120 32376 27126 32428
rect 28258 32308 28264 32360
rect 28316 32308 28322 32360
rect 23900 32252 25084 32280
rect 23900 32240 23906 32252
rect 7248 32184 7880 32212
rect 11793 32215 11851 32221
rect 7248 32172 7254 32184
rect 11793 32181 11805 32215
rect 11839 32212 11851 32215
rect 12250 32212 12256 32224
rect 11839 32184 12256 32212
rect 11839 32181 11851 32184
rect 11793 32175 11851 32181
rect 12250 32172 12256 32184
rect 12308 32172 12314 32224
rect 18782 32172 18788 32224
rect 18840 32212 18846 32224
rect 19061 32215 19119 32221
rect 19061 32212 19073 32215
rect 18840 32184 19073 32212
rect 18840 32172 18846 32184
rect 19061 32181 19073 32184
rect 19107 32181 19119 32215
rect 19061 32175 19119 32181
rect 22186 32172 22192 32224
rect 22244 32212 22250 32224
rect 22741 32215 22799 32221
rect 22741 32212 22753 32215
rect 22244 32184 22753 32212
rect 22244 32172 22250 32184
rect 22741 32181 22753 32184
rect 22787 32181 22799 32215
rect 22741 32175 22799 32181
rect 23106 32172 23112 32224
rect 23164 32172 23170 32224
rect 23569 32215 23627 32221
rect 23569 32181 23581 32215
rect 23615 32212 23627 32215
rect 25038 32212 25044 32224
rect 23615 32184 25044 32212
rect 23615 32181 23627 32184
rect 23569 32175 23627 32181
rect 25038 32172 25044 32184
rect 25096 32172 25102 32224
rect 25130 32172 25136 32224
rect 25188 32212 25194 32224
rect 25593 32215 25651 32221
rect 25593 32212 25605 32215
rect 25188 32184 25605 32212
rect 25188 32172 25194 32184
rect 25593 32181 25605 32184
rect 25639 32212 25651 32215
rect 25774 32212 25780 32224
rect 25639 32184 25780 32212
rect 25639 32181 25651 32184
rect 25593 32175 25651 32181
rect 25774 32172 25780 32184
rect 25832 32172 25838 32224
rect 1104 32122 28888 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 28888 32122
rect 1104 32048 28888 32070
rect 5994 31968 6000 32020
rect 6052 32008 6058 32020
rect 7009 32011 7067 32017
rect 7009 32008 7021 32011
rect 6052 31980 7021 32008
rect 6052 31968 6058 31980
rect 7009 31977 7021 31980
rect 7055 31977 7067 32011
rect 7009 31971 7067 31977
rect 7926 31968 7932 32020
rect 7984 31968 7990 32020
rect 12710 31968 12716 32020
rect 12768 31968 12774 32020
rect 15286 31968 15292 32020
rect 15344 32008 15350 32020
rect 15381 32011 15439 32017
rect 15381 32008 15393 32011
rect 15344 31980 15393 32008
rect 15344 31968 15350 31980
rect 15381 31977 15393 31980
rect 15427 31977 15439 32011
rect 15381 31971 15439 31977
rect 16669 32011 16727 32017
rect 16669 31977 16681 32011
rect 16715 32008 16727 32011
rect 17034 32008 17040 32020
rect 16715 31980 17040 32008
rect 16715 31977 16727 31980
rect 16669 31971 16727 31977
rect 17034 31968 17040 31980
rect 17092 31968 17098 32020
rect 18598 31968 18604 32020
rect 18656 31968 18662 32020
rect 19889 32011 19947 32017
rect 19889 31977 19901 32011
rect 19935 32008 19947 32011
rect 21082 32008 21088 32020
rect 19935 31980 21088 32008
rect 19935 31977 19947 31980
rect 19889 31971 19947 31977
rect 21082 31968 21088 31980
rect 21140 31968 21146 32020
rect 21174 31968 21180 32020
rect 21232 31968 21238 32020
rect 22281 32011 22339 32017
rect 22066 31980 22232 32008
rect 6733 31943 6791 31949
rect 6733 31909 6745 31943
rect 6779 31940 6791 31943
rect 22066 31940 22094 31980
rect 6779 31912 6914 31940
rect 6779 31909 6791 31912
rect 6733 31903 6791 31909
rect 6886 31872 6914 31912
rect 21008 31912 22094 31940
rect 22204 31940 22232 31980
rect 22281 31977 22293 32011
rect 22327 32008 22339 32011
rect 23750 32008 23756 32020
rect 22327 31980 23756 32008
rect 22327 31977 22339 31980
rect 22281 31971 22339 31977
rect 23750 31968 23756 31980
rect 23808 31968 23814 32020
rect 22204 31912 22968 31940
rect 7561 31875 7619 31881
rect 7561 31872 7573 31875
rect 6886 31844 7573 31872
rect 7561 31841 7573 31844
rect 7607 31841 7619 31875
rect 8573 31875 8631 31881
rect 8573 31872 8585 31875
rect 7561 31835 7619 31841
rect 8128 31844 8585 31872
rect 5353 31807 5411 31813
rect 5353 31773 5365 31807
rect 5399 31804 5411 31807
rect 7190 31804 7196 31816
rect 5399 31776 7196 31804
rect 5399 31773 5411 31776
rect 5353 31767 5411 31773
rect 7190 31764 7196 31776
rect 7248 31764 7254 31816
rect 8128 31813 8156 31844
rect 8573 31841 8585 31844
rect 8619 31841 8631 31875
rect 8573 31835 8631 31841
rect 16390 31832 16396 31884
rect 16448 31872 16454 31884
rect 16761 31875 16819 31881
rect 16761 31872 16773 31875
rect 16448 31844 16773 31872
rect 16448 31832 16454 31844
rect 16761 31841 16773 31844
rect 16807 31841 16819 31875
rect 16761 31835 16819 31841
rect 19242 31832 19248 31884
rect 19300 31872 19306 31884
rect 19521 31875 19579 31881
rect 19521 31872 19533 31875
rect 19300 31844 19533 31872
rect 19300 31832 19306 31844
rect 19521 31841 19533 31844
rect 19567 31841 19579 31875
rect 19521 31835 19579 31841
rect 19702 31832 19708 31884
rect 19760 31832 19766 31884
rect 21008 31881 21036 31912
rect 20625 31875 20683 31881
rect 20625 31841 20637 31875
rect 20671 31872 20683 31875
rect 20993 31875 21051 31881
rect 20993 31872 21005 31875
rect 20671 31844 21005 31872
rect 20671 31841 20683 31844
rect 20625 31835 20683 31841
rect 20993 31841 21005 31844
rect 21039 31841 21051 31875
rect 20993 31835 21051 31841
rect 21821 31875 21879 31881
rect 21821 31841 21833 31875
rect 21867 31872 21879 31875
rect 22186 31872 22192 31884
rect 21867 31844 22192 31872
rect 21867 31841 21879 31844
rect 21821 31835 21879 31841
rect 22186 31832 22192 31844
rect 22244 31832 22250 31884
rect 22940 31881 22968 31912
rect 22925 31875 22983 31881
rect 22925 31841 22937 31875
rect 22971 31841 22983 31875
rect 22925 31835 22983 31841
rect 8113 31807 8171 31813
rect 8113 31773 8125 31807
rect 8159 31773 8171 31807
rect 8113 31767 8171 31773
rect 5626 31745 5632 31748
rect 5620 31736 5632 31745
rect 5587 31708 5632 31736
rect 5620 31699 5632 31708
rect 5626 31696 5632 31699
rect 5684 31696 5690 31748
rect 6638 31696 6644 31748
rect 6696 31736 6702 31748
rect 8128 31736 8156 31767
rect 8294 31764 8300 31816
rect 8352 31764 8358 31816
rect 12158 31764 12164 31816
rect 12216 31804 12222 31816
rect 12621 31807 12679 31813
rect 12621 31804 12633 31807
rect 12216 31776 12633 31804
rect 12216 31764 12222 31776
rect 12621 31773 12633 31776
rect 12667 31773 12679 31807
rect 12621 31767 12679 31773
rect 12802 31764 12808 31816
rect 12860 31764 12866 31816
rect 16025 31807 16083 31813
rect 16025 31773 16037 31807
rect 16071 31804 16083 31807
rect 16301 31807 16359 31813
rect 16301 31804 16313 31807
rect 16071 31776 16313 31804
rect 16071 31773 16083 31776
rect 16025 31767 16083 31773
rect 16301 31773 16313 31776
rect 16347 31773 16359 31807
rect 16301 31767 16359 31773
rect 16482 31764 16488 31816
rect 16540 31764 16546 31816
rect 18782 31764 18788 31816
rect 18840 31764 18846 31816
rect 18874 31764 18880 31816
rect 18932 31804 18938 31816
rect 18932 31776 19196 31804
rect 18932 31764 18938 31776
rect 6696 31708 8156 31736
rect 6696 31696 6702 31708
rect 18598 31696 18604 31748
rect 18656 31696 18662 31748
rect 19168 31736 19196 31776
rect 19426 31764 19432 31816
rect 19484 31764 19490 31816
rect 19610 31764 19616 31816
rect 19668 31764 19674 31816
rect 20533 31807 20591 31813
rect 20533 31804 20545 31807
rect 19812 31776 20545 31804
rect 19812 31754 19840 31776
rect 20533 31773 20545 31776
rect 20579 31804 20591 31807
rect 20717 31807 20775 31813
rect 20579 31776 20668 31804
rect 20579 31773 20591 31776
rect 20533 31767 20591 31773
rect 19720 31736 19840 31754
rect 19168 31726 19840 31736
rect 20640 31736 20668 31776
rect 20717 31773 20729 31807
rect 20763 31804 20775 31807
rect 20763 31776 20944 31804
rect 20763 31773 20775 31776
rect 20717 31767 20775 31773
rect 20806 31736 20812 31748
rect 19168 31708 19748 31726
rect 20640 31708 20812 31736
rect 20806 31696 20812 31708
rect 20864 31696 20870 31748
rect 20916 31668 20944 31776
rect 21082 31764 21088 31816
rect 21140 31804 21146 31816
rect 21450 31804 21456 31816
rect 21140 31776 21456 31804
rect 21140 31764 21146 31776
rect 21450 31764 21456 31776
rect 21508 31764 21514 31816
rect 21913 31807 21971 31813
rect 21913 31804 21925 31807
rect 21891 31776 21925 31804
rect 21913 31773 21925 31776
rect 21959 31773 21971 31807
rect 21913 31767 21971 31773
rect 21174 31696 21180 31748
rect 21232 31736 21238 31748
rect 21361 31739 21419 31745
rect 21361 31736 21373 31739
rect 21232 31708 21373 31736
rect 21232 31696 21238 31708
rect 21361 31705 21373 31708
rect 21407 31736 21419 31739
rect 21928 31736 21956 31767
rect 22002 31764 22008 31816
rect 22060 31764 22066 31816
rect 22094 31764 22100 31816
rect 22152 31764 22158 31816
rect 22557 31807 22615 31813
rect 22557 31804 22569 31807
rect 22204 31776 22569 31804
rect 22204 31736 22232 31776
rect 22557 31773 22569 31776
rect 22603 31773 22615 31807
rect 22557 31767 22615 31773
rect 22738 31764 22744 31816
rect 22796 31764 22802 31816
rect 23566 31764 23572 31816
rect 23624 31804 23630 31816
rect 24121 31807 24179 31813
rect 24121 31804 24133 31807
rect 23624 31776 24133 31804
rect 23624 31764 23630 31776
rect 24121 31773 24133 31776
rect 24167 31804 24179 31807
rect 24578 31804 24584 31816
rect 24167 31776 24584 31804
rect 24167 31773 24179 31776
rect 24121 31767 24179 31773
rect 24578 31764 24584 31776
rect 24636 31764 24642 31816
rect 28442 31764 28448 31816
rect 28500 31764 28506 31816
rect 21407 31708 22232 31736
rect 21407 31705 21419 31708
rect 21361 31699 21419 31705
rect 22094 31668 22100 31680
rect 20916 31640 22100 31668
rect 22094 31628 22100 31640
rect 22152 31628 22158 31680
rect 1104 31578 28888 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 28888 31578
rect 1104 31504 28888 31526
rect 7837 31467 7895 31473
rect 7837 31433 7849 31467
rect 7883 31464 7895 31467
rect 8294 31464 8300 31476
rect 7883 31436 8300 31464
rect 7883 31433 7895 31436
rect 7837 31427 7895 31433
rect 8294 31424 8300 31436
rect 8352 31424 8358 31476
rect 22281 31467 22339 31473
rect 22281 31433 22293 31467
rect 22327 31464 22339 31467
rect 22738 31464 22744 31476
rect 22327 31436 22744 31464
rect 22327 31433 22339 31436
rect 22281 31427 22339 31433
rect 22738 31424 22744 31436
rect 22796 31424 22802 31476
rect 20806 31356 20812 31408
rect 20864 31396 20870 31408
rect 21910 31396 21916 31408
rect 20864 31368 21916 31396
rect 20864 31356 20870 31368
rect 21910 31356 21916 31368
rect 21968 31356 21974 31408
rect 22094 31356 22100 31408
rect 22152 31356 22158 31408
rect 5902 31288 5908 31340
rect 5960 31328 5966 31340
rect 6457 31331 6515 31337
rect 6457 31328 6469 31331
rect 5960 31300 6469 31328
rect 5960 31288 5966 31300
rect 6457 31297 6469 31300
rect 6503 31297 6515 31331
rect 6457 31291 6515 31297
rect 6638 31288 6644 31340
rect 6696 31288 6702 31340
rect 6822 31288 6828 31340
rect 6880 31328 6886 31340
rect 7193 31331 7251 31337
rect 7193 31328 7205 31331
rect 6880 31300 7205 31328
rect 6880 31288 6886 31300
rect 7193 31297 7205 31300
rect 7239 31297 7251 31331
rect 7193 31291 7251 31297
rect 21174 31288 21180 31340
rect 21232 31288 21238 31340
rect 21269 31263 21327 31269
rect 21269 31229 21281 31263
rect 21315 31260 21327 31263
rect 21450 31260 21456 31272
rect 21315 31232 21456 31260
rect 21315 31229 21327 31232
rect 21269 31223 21327 31229
rect 21450 31220 21456 31232
rect 21508 31260 21514 31272
rect 22002 31260 22008 31272
rect 21508 31232 22008 31260
rect 21508 31220 21514 31232
rect 22002 31220 22008 31232
rect 22060 31220 22066 31272
rect 21542 31152 21548 31204
rect 21600 31152 21606 31204
rect 6822 31084 6828 31136
rect 6880 31084 6886 31136
rect 1104 31034 28888 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 28888 31034
rect 1104 30960 28888 30982
rect 5537 30923 5595 30929
rect 5537 30889 5549 30923
rect 5583 30920 5595 30923
rect 6730 30920 6736 30932
rect 5583 30892 6736 30920
rect 5583 30889 5595 30892
rect 5537 30883 5595 30889
rect 6730 30880 6736 30892
rect 6788 30880 6794 30932
rect 18598 30880 18604 30932
rect 18656 30880 18662 30932
rect 19610 30784 19616 30796
rect 18800 30756 19616 30784
rect 6661 30719 6719 30725
rect 6661 30685 6673 30719
rect 6707 30716 6719 30719
rect 6822 30716 6828 30728
rect 6707 30688 6828 30716
rect 6707 30685 6719 30688
rect 6661 30679 6719 30685
rect 6822 30676 6828 30688
rect 6880 30676 6886 30728
rect 6917 30719 6975 30725
rect 6917 30685 6929 30719
rect 6963 30716 6975 30719
rect 7190 30716 7196 30728
rect 6963 30688 7196 30716
rect 6963 30685 6975 30688
rect 6917 30679 6975 30685
rect 7190 30676 7196 30688
rect 7248 30676 7254 30728
rect 18800 30725 18828 30756
rect 19610 30744 19616 30756
rect 19668 30744 19674 30796
rect 18785 30719 18843 30725
rect 18785 30685 18797 30719
rect 18831 30685 18843 30719
rect 18785 30679 18843 30685
rect 18877 30719 18935 30725
rect 18877 30685 18889 30719
rect 18923 30716 18935 30719
rect 19242 30716 19248 30728
rect 18923 30688 19248 30716
rect 18923 30685 18935 30688
rect 18877 30679 18935 30685
rect 17678 30608 17684 30660
rect 17736 30648 17742 30660
rect 18892 30648 18920 30679
rect 19242 30676 19248 30688
rect 19300 30676 19306 30728
rect 17736 30620 18920 30648
rect 17736 30608 17742 30620
rect 6638 30540 6644 30592
rect 6696 30580 6702 30592
rect 7285 30583 7343 30589
rect 7285 30580 7297 30583
rect 6696 30552 7297 30580
rect 6696 30540 6702 30552
rect 7285 30549 7297 30552
rect 7331 30580 7343 30583
rect 8478 30580 8484 30592
rect 7331 30552 8484 30580
rect 7331 30549 7343 30552
rect 7285 30543 7343 30549
rect 8478 30540 8484 30552
rect 8536 30540 8542 30592
rect 17589 30583 17647 30589
rect 17589 30549 17601 30583
rect 17635 30580 17647 30583
rect 17770 30580 17776 30592
rect 17635 30552 17776 30580
rect 17635 30549 17647 30552
rect 17589 30543 17647 30549
rect 17770 30540 17776 30552
rect 17828 30540 17834 30592
rect 1104 30490 28888 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 28888 30490
rect 1104 30416 28888 30438
rect 17865 30311 17923 30317
rect 17865 30277 17877 30311
rect 17911 30308 17923 30311
rect 18233 30311 18291 30317
rect 18233 30308 18245 30311
rect 17911 30280 18245 30308
rect 17911 30277 17923 30280
rect 17865 30271 17923 30277
rect 18233 30277 18245 30280
rect 18279 30277 18291 30311
rect 18233 30271 18291 30277
rect 18417 30311 18475 30317
rect 18417 30277 18429 30311
rect 18463 30308 18475 30311
rect 18598 30308 18604 30320
rect 18463 30280 18604 30308
rect 18463 30277 18475 30280
rect 18417 30271 18475 30277
rect 18598 30268 18604 30280
rect 18656 30268 18662 30320
rect 24210 30268 24216 30320
rect 24268 30268 24274 30320
rect 1302 30200 1308 30252
rect 1360 30240 1366 30252
rect 1489 30243 1547 30249
rect 1489 30240 1501 30243
rect 1360 30212 1501 30240
rect 1360 30200 1366 30212
rect 1489 30209 1501 30212
rect 1535 30240 1547 30243
rect 1949 30243 2007 30249
rect 1949 30240 1961 30243
rect 1535 30212 1961 30240
rect 1535 30209 1547 30212
rect 1489 30203 1547 30209
rect 1949 30209 1961 30212
rect 1995 30209 2007 30243
rect 1949 30203 2007 30209
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30209 17371 30243
rect 17313 30203 17371 30209
rect 17497 30243 17555 30249
rect 17497 30209 17509 30243
rect 17543 30209 17555 30243
rect 17497 30203 17555 30209
rect 9030 30132 9036 30184
rect 9088 30172 9094 30184
rect 9953 30175 10011 30181
rect 9953 30172 9965 30175
rect 9088 30144 9965 30172
rect 9088 30132 9094 30144
rect 9953 30141 9965 30144
rect 9999 30141 10011 30175
rect 9953 30135 10011 30141
rect 17328 30116 17356 30203
rect 17512 30172 17540 30203
rect 17678 30200 17684 30252
rect 17736 30240 17742 30252
rect 17773 30243 17831 30249
rect 17773 30240 17785 30243
rect 17736 30212 17785 30240
rect 17736 30200 17742 30212
rect 17773 30209 17785 30212
rect 17819 30209 17831 30243
rect 17773 30203 17831 30209
rect 17957 30243 18015 30249
rect 17957 30209 17969 30243
rect 18003 30240 18015 30243
rect 19610 30240 19616 30252
rect 18003 30212 19616 30240
rect 18003 30209 18015 30212
rect 17957 30203 18015 30209
rect 19610 30200 19616 30212
rect 19668 30200 19674 30252
rect 23750 30200 23756 30252
rect 23808 30200 23814 30252
rect 23842 30200 23848 30252
rect 23900 30200 23906 30252
rect 24029 30243 24087 30249
rect 24029 30209 24041 30243
rect 24075 30240 24087 30243
rect 24118 30240 24124 30252
rect 24075 30212 24124 30240
rect 24075 30209 24087 30212
rect 24029 30203 24087 30209
rect 24118 30200 24124 30212
rect 24176 30200 24182 30252
rect 18877 30175 18935 30181
rect 18877 30172 18889 30175
rect 17512 30144 18889 30172
rect 18877 30141 18889 30144
rect 18923 30141 18935 30175
rect 18877 30135 18935 30141
rect 19334 30132 19340 30184
rect 19392 30172 19398 30184
rect 19429 30175 19487 30181
rect 19429 30172 19441 30175
rect 19392 30144 19441 30172
rect 19392 30132 19398 30144
rect 19429 30141 19441 30144
rect 19475 30141 19487 30175
rect 19429 30135 19487 30141
rect 17310 30064 17316 30116
rect 17368 30104 17374 30116
rect 17770 30104 17776 30116
rect 17368 30076 17776 30104
rect 17368 30064 17374 30076
rect 17770 30064 17776 30076
rect 17828 30104 17834 30116
rect 20622 30104 20628 30116
rect 17828 30076 20628 30104
rect 17828 30064 17834 30076
rect 20622 30064 20628 30076
rect 20680 30064 20686 30116
rect 1670 29996 1676 30048
rect 1728 29996 1734 30048
rect 8478 29996 8484 30048
rect 8536 30036 8542 30048
rect 8757 30039 8815 30045
rect 8757 30036 8769 30039
rect 8536 30008 8769 30036
rect 8536 29996 8542 30008
rect 8757 30005 8769 30008
rect 8803 30005 8815 30039
rect 8757 29999 8815 30005
rect 9398 29996 9404 30048
rect 9456 29996 9462 30048
rect 17494 29996 17500 30048
rect 17552 29996 17558 30048
rect 18598 29996 18604 30048
rect 18656 29996 18662 30048
rect 1104 29946 28888 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 28888 29946
rect 1104 29872 28888 29894
rect 10689 29835 10747 29841
rect 10689 29832 10701 29835
rect 8312 29804 10701 29832
rect 8312 29705 8340 29804
rect 10689 29801 10701 29804
rect 10735 29801 10747 29835
rect 10689 29795 10747 29801
rect 15102 29792 15108 29844
rect 15160 29832 15166 29844
rect 15473 29835 15531 29841
rect 15473 29832 15485 29835
rect 15160 29804 15485 29832
rect 15160 29792 15166 29804
rect 15473 29801 15485 29804
rect 15519 29832 15531 29835
rect 17310 29832 17316 29844
rect 15519 29804 17316 29832
rect 15519 29801 15531 29804
rect 15473 29795 15531 29801
rect 17310 29792 17316 29804
rect 17368 29792 17374 29844
rect 18782 29792 18788 29844
rect 18840 29832 18846 29844
rect 18969 29835 19027 29841
rect 18969 29832 18981 29835
rect 18840 29804 18981 29832
rect 18840 29792 18846 29804
rect 18969 29801 18981 29804
rect 19015 29801 19027 29835
rect 18969 29795 19027 29801
rect 19334 29792 19340 29844
rect 19392 29792 19398 29844
rect 24578 29792 24584 29844
rect 24636 29792 24642 29844
rect 9030 29724 9036 29776
rect 9088 29724 9094 29776
rect 8297 29699 8355 29705
rect 8297 29665 8309 29699
rect 8343 29665 8355 29699
rect 8297 29659 8355 29665
rect 10502 29656 10508 29708
rect 10560 29696 10566 29708
rect 11241 29699 11299 29705
rect 11241 29696 11253 29699
rect 10560 29668 11253 29696
rect 10560 29656 10566 29668
rect 11241 29665 11253 29668
rect 11287 29665 11299 29699
rect 11241 29659 11299 29665
rect 17586 29656 17592 29708
rect 17644 29656 17650 29708
rect 18598 29656 18604 29708
rect 18656 29696 18662 29708
rect 19797 29699 19855 29705
rect 19797 29696 19809 29699
rect 18656 29668 19809 29696
rect 18656 29656 18662 29668
rect 19797 29665 19809 29668
rect 19843 29665 19855 29699
rect 19797 29659 19855 29665
rect 19886 29656 19892 29708
rect 19944 29656 19950 29708
rect 21910 29656 21916 29708
rect 21968 29696 21974 29708
rect 21968 29668 23980 29696
rect 21968 29656 21974 29668
rect 842 29588 848 29640
rect 900 29628 906 29640
rect 1489 29631 1547 29637
rect 1489 29628 1501 29631
rect 900 29600 1501 29628
rect 900 29588 906 29600
rect 1489 29597 1501 29600
rect 1535 29597 1547 29631
rect 1489 29591 1547 29597
rect 8478 29588 8484 29640
rect 8536 29588 8542 29640
rect 10318 29588 10324 29640
rect 10376 29628 10382 29640
rect 10413 29631 10471 29637
rect 10413 29628 10425 29631
rect 10376 29600 10425 29628
rect 10376 29588 10382 29600
rect 10413 29597 10425 29600
rect 10459 29597 10471 29631
rect 10413 29591 10471 29597
rect 17494 29588 17500 29640
rect 17552 29628 17558 29640
rect 23952 29637 23980 29668
rect 17845 29631 17903 29637
rect 17845 29628 17857 29631
rect 17552 29600 17857 29628
rect 17552 29588 17558 29600
rect 17845 29597 17857 29600
rect 17891 29597 17903 29631
rect 17845 29591 17903 29597
rect 23845 29631 23903 29637
rect 23845 29597 23857 29631
rect 23891 29597 23903 29631
rect 23845 29591 23903 29597
rect 23937 29631 23995 29637
rect 23937 29597 23949 29631
rect 23983 29597 23995 29631
rect 23937 29591 23995 29597
rect 8665 29563 8723 29569
rect 8665 29529 8677 29563
rect 8711 29560 8723 29563
rect 10146 29563 10204 29569
rect 10146 29560 10158 29563
rect 8711 29532 10158 29560
rect 8711 29529 8723 29532
rect 8665 29523 8723 29529
rect 10146 29529 10158 29532
rect 10192 29529 10204 29563
rect 23860 29560 23888 29591
rect 24946 29560 24952 29572
rect 23860 29532 24952 29560
rect 10146 29523 10204 29529
rect 24946 29520 24952 29532
rect 25004 29520 25010 29572
rect 19426 29452 19432 29504
rect 19484 29492 19490 29504
rect 19705 29495 19763 29501
rect 19705 29492 19717 29495
rect 19484 29464 19717 29492
rect 19484 29452 19490 29464
rect 19705 29461 19717 29464
rect 19751 29461 19763 29495
rect 19705 29455 19763 29461
rect 24118 29452 24124 29504
rect 24176 29452 24182 29504
rect 1104 29402 28888 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 28888 29402
rect 1104 29328 28888 29350
rect 9766 29248 9772 29300
rect 9824 29288 9830 29300
rect 9861 29291 9919 29297
rect 9861 29288 9873 29291
rect 9824 29260 9873 29288
rect 9824 29248 9830 29260
rect 9861 29257 9873 29260
rect 9907 29288 9919 29291
rect 10502 29288 10508 29300
rect 9907 29260 10508 29288
rect 9907 29257 9919 29260
rect 9861 29251 9919 29257
rect 10502 29248 10508 29260
rect 10560 29248 10566 29300
rect 18325 29291 18383 29297
rect 18325 29257 18337 29291
rect 18371 29288 18383 29291
rect 19610 29288 19616 29300
rect 18371 29260 19616 29288
rect 18371 29257 18383 29260
rect 18325 29251 18383 29257
rect 19610 29248 19616 29260
rect 19668 29248 19674 29300
rect 24946 29288 24952 29300
rect 23124 29260 24952 29288
rect 8294 29180 8300 29232
rect 8352 29220 8358 29232
rect 8352 29192 9168 29220
rect 8352 29180 8358 29192
rect 1670 29112 1676 29164
rect 1728 29152 1734 29164
rect 3789 29155 3847 29161
rect 3789 29152 3801 29155
rect 1728 29124 3801 29152
rect 1728 29112 1734 29124
rect 3789 29121 3801 29124
rect 3835 29121 3847 29155
rect 3789 29115 3847 29121
rect 7653 29155 7711 29161
rect 7653 29121 7665 29155
rect 7699 29152 7711 29155
rect 8113 29155 8171 29161
rect 8113 29152 8125 29155
rect 7699 29124 8125 29152
rect 7699 29121 7711 29124
rect 7653 29115 7711 29121
rect 8113 29121 8125 29124
rect 8159 29152 8171 29155
rect 8478 29152 8484 29164
rect 8159 29124 8484 29152
rect 8159 29121 8171 29124
rect 8113 29115 8171 29121
rect 3605 29087 3663 29093
rect 3605 29053 3617 29087
rect 3651 29084 3663 29087
rect 4341 29087 4399 29093
rect 4341 29084 4353 29087
rect 3651 29056 4353 29084
rect 3651 29053 3663 29056
rect 3605 29047 3663 29053
rect 4341 29053 4353 29056
rect 4387 29084 4399 29087
rect 7668 29084 7696 29115
rect 8478 29112 8484 29124
rect 8536 29112 8542 29164
rect 9140 29161 9168 29192
rect 10870 29180 10876 29232
rect 10928 29220 10934 29232
rect 10974 29223 11032 29229
rect 10974 29220 10986 29223
rect 10928 29192 10986 29220
rect 10928 29180 10934 29192
rect 10974 29189 10986 29192
rect 11020 29189 11032 29223
rect 10974 29183 11032 29189
rect 12621 29223 12679 29229
rect 12621 29189 12633 29223
rect 12667 29220 12679 29223
rect 12894 29220 12900 29232
rect 12667 29192 12900 29220
rect 12667 29189 12679 29192
rect 12621 29183 12679 29189
rect 12894 29180 12900 29192
rect 12952 29220 12958 29232
rect 13538 29220 13544 29232
rect 12952 29192 13544 29220
rect 12952 29180 12958 29192
rect 13538 29180 13544 29192
rect 13596 29180 13602 29232
rect 14369 29223 14427 29229
rect 14369 29220 14381 29223
rect 13740 29192 14381 29220
rect 9125 29155 9183 29161
rect 9125 29121 9137 29155
rect 9171 29121 9183 29155
rect 9125 29115 9183 29121
rect 12986 29112 12992 29164
rect 13044 29152 13050 29164
rect 13265 29155 13323 29161
rect 13265 29152 13277 29155
rect 13044 29124 13277 29152
rect 13044 29112 13050 29124
rect 13265 29121 13277 29124
rect 13311 29121 13323 29155
rect 13265 29115 13323 29121
rect 13630 29112 13636 29164
rect 13688 29152 13694 29164
rect 13740 29161 13768 29192
rect 14369 29189 14381 29192
rect 14415 29189 14427 29223
rect 18138 29220 18144 29232
rect 14369 29183 14427 29189
rect 16546 29192 18144 29220
rect 13725 29155 13783 29161
rect 13725 29152 13737 29155
rect 13688 29124 13737 29152
rect 13688 29112 13694 29124
rect 13725 29121 13737 29124
rect 13771 29121 13783 29155
rect 13725 29115 13783 29121
rect 13814 29112 13820 29164
rect 13872 29152 13878 29164
rect 13909 29155 13967 29161
rect 13909 29152 13921 29155
rect 13872 29124 13921 29152
rect 13872 29112 13878 29124
rect 13909 29121 13921 29124
rect 13955 29152 13967 29155
rect 14185 29155 14243 29161
rect 14185 29152 14197 29155
rect 13955 29124 14197 29152
rect 13955 29121 13967 29124
rect 13909 29115 13967 29121
rect 14185 29121 14197 29124
rect 14231 29121 14243 29155
rect 14185 29115 14243 29121
rect 15102 29112 15108 29164
rect 15160 29112 15166 29164
rect 15286 29112 15292 29164
rect 15344 29112 15350 29164
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29152 15899 29155
rect 16390 29152 16396 29164
rect 15887 29124 16396 29152
rect 15887 29121 15899 29124
rect 15841 29115 15899 29121
rect 16390 29112 16396 29124
rect 16448 29152 16454 29164
rect 16546 29152 16574 29192
rect 18138 29180 18144 29192
rect 18196 29180 18202 29232
rect 21910 29220 21916 29232
rect 18616 29192 21916 29220
rect 16448 29124 16574 29152
rect 16448 29112 16454 29124
rect 16758 29112 16764 29164
rect 16816 29112 16822 29164
rect 16942 29112 16948 29164
rect 17000 29112 17006 29164
rect 4387 29056 7696 29084
rect 7929 29087 7987 29093
rect 4387 29053 4399 29056
rect 4341 29047 4399 29053
rect 7929 29053 7941 29087
rect 7975 29084 7987 29087
rect 8573 29087 8631 29093
rect 8573 29084 8585 29087
rect 7975 29056 8585 29084
rect 7975 29053 7987 29056
rect 7929 29047 7987 29053
rect 8573 29053 8585 29056
rect 8619 29053 8631 29087
rect 8573 29047 8631 29053
rect 11241 29087 11299 29093
rect 11241 29053 11253 29087
rect 11287 29053 11299 29087
rect 11241 29047 11299 29053
rect 3973 29019 4031 29025
rect 3973 28985 3985 29019
rect 4019 29016 4031 29019
rect 4798 29016 4804 29028
rect 4019 28988 4804 29016
rect 4019 28985 4031 28988
rect 3973 28979 4031 28985
rect 4798 28976 4804 28988
rect 4856 28976 4862 29028
rect 8297 29019 8355 29025
rect 8297 28985 8309 29019
rect 8343 29016 8355 29019
rect 10042 29016 10048 29028
rect 8343 28988 10048 29016
rect 8343 28985 8355 28988
rect 8297 28979 8355 28985
rect 10042 28976 10048 28988
rect 10100 28976 10106 29028
rect 9858 28908 9864 28960
rect 9916 28948 9922 28960
rect 10318 28948 10324 28960
rect 9916 28920 10324 28948
rect 9916 28908 9922 28920
rect 10318 28908 10324 28920
rect 10376 28948 10382 28960
rect 10962 28948 10968 28960
rect 10376 28920 10968 28948
rect 10376 28908 10382 28920
rect 10962 28908 10968 28920
rect 11020 28948 11026 28960
rect 11256 28948 11284 29047
rect 11330 29044 11336 29096
rect 11388 29084 11394 29096
rect 12161 29087 12219 29093
rect 12161 29084 12173 29087
rect 11388 29056 12173 29084
rect 11388 29044 11394 29056
rect 12161 29053 12173 29056
rect 12207 29053 12219 29087
rect 12161 29047 12219 29053
rect 15194 29044 15200 29096
rect 15252 29044 15258 29096
rect 15933 29087 15991 29093
rect 15933 29053 15945 29087
rect 15979 29084 15991 29087
rect 16853 29087 16911 29093
rect 16853 29084 16865 29087
rect 15979 29056 16865 29084
rect 15979 29053 15991 29056
rect 15933 29047 15991 29053
rect 16853 29053 16865 29056
rect 16899 29053 16911 29087
rect 16853 29047 16911 29053
rect 17954 29044 17960 29096
rect 18012 29084 18018 29096
rect 18616 29093 18644 29192
rect 21910 29180 21916 29192
rect 21968 29220 21974 29232
rect 23124 29229 23152 29260
rect 24946 29248 24952 29260
rect 25004 29248 25010 29300
rect 26697 29291 26755 29297
rect 26697 29257 26709 29291
rect 26743 29288 26755 29291
rect 27062 29288 27068 29300
rect 26743 29260 27068 29288
rect 26743 29257 26755 29260
rect 26697 29251 26755 29257
rect 27062 29248 27068 29260
rect 27120 29248 27126 29300
rect 22925 29223 22983 29229
rect 22925 29220 22937 29223
rect 21968 29192 22937 29220
rect 21968 29180 21974 29192
rect 22925 29189 22937 29192
rect 22971 29189 22983 29223
rect 22925 29183 22983 29189
rect 23109 29223 23167 29229
rect 23109 29189 23121 29223
rect 23155 29189 23167 29223
rect 23109 29183 23167 29189
rect 24118 29180 24124 29232
rect 24176 29220 24182 29232
rect 24857 29223 24915 29229
rect 24857 29220 24869 29223
rect 24176 29192 24869 29220
rect 24176 29180 24182 29192
rect 24857 29189 24869 29192
rect 24903 29189 24915 29223
rect 24857 29183 24915 29189
rect 18693 29155 18751 29161
rect 18693 29121 18705 29155
rect 18739 29121 18751 29155
rect 18693 29115 18751 29121
rect 18601 29087 18659 29093
rect 18601 29084 18613 29087
rect 18012 29056 18613 29084
rect 18012 29044 18018 29056
rect 18601 29053 18613 29056
rect 18647 29053 18659 29087
rect 18708 29084 18736 29115
rect 18782 29112 18788 29164
rect 18840 29152 18846 29164
rect 19153 29155 19211 29161
rect 19153 29152 19165 29155
rect 18840 29124 19165 29152
rect 18840 29112 18846 29124
rect 19153 29121 19165 29124
rect 19199 29121 19211 29155
rect 19153 29115 19211 29121
rect 23753 29155 23811 29161
rect 23753 29121 23765 29155
rect 23799 29152 23811 29155
rect 23799 29124 24440 29152
rect 23799 29121 23811 29124
rect 23753 29115 23811 29121
rect 19426 29084 19432 29096
rect 18708 29056 19432 29084
rect 18601 29047 18659 29053
rect 19426 29044 19432 29056
rect 19484 29044 19490 29096
rect 23658 29044 23664 29096
rect 23716 29044 23722 29096
rect 24412 29093 24440 29124
rect 25314 29112 25320 29164
rect 25372 29112 25378 29164
rect 25584 29155 25642 29161
rect 25584 29121 25596 29155
rect 25630 29152 25642 29155
rect 26050 29152 26056 29164
rect 25630 29124 26056 29152
rect 25630 29121 25642 29124
rect 25584 29115 25642 29121
rect 26050 29112 26056 29124
rect 26108 29112 26114 29164
rect 24397 29087 24455 29093
rect 24397 29053 24409 29087
rect 24443 29053 24455 29087
rect 24397 29047 24455 29053
rect 13817 29019 13875 29025
rect 13817 28985 13829 29019
rect 13863 29016 13875 29019
rect 14366 29016 14372 29028
rect 13863 28988 14372 29016
rect 13863 28985 13875 28988
rect 13817 28979 13875 28985
rect 14366 28976 14372 28988
rect 14424 28976 14430 29028
rect 14553 29019 14611 29025
rect 14553 28985 14565 29019
rect 14599 29016 14611 29019
rect 14734 29016 14740 29028
rect 14599 28988 14740 29016
rect 14599 28985 14611 28988
rect 14553 28979 14611 28985
rect 14734 28976 14740 28988
rect 14792 28976 14798 29028
rect 16209 29019 16267 29025
rect 16209 28985 16221 29019
rect 16255 29016 16267 29019
rect 16758 29016 16764 29028
rect 16255 28988 16764 29016
rect 16255 28985 16267 28988
rect 16209 28979 16267 28985
rect 16758 28976 16764 28988
rect 16816 28976 16822 29028
rect 19886 29016 19892 29028
rect 19444 28988 19892 29016
rect 11020 28920 11284 28948
rect 11020 28908 11026 28920
rect 11422 28908 11428 28960
rect 11480 28948 11486 28960
rect 11609 28951 11667 28957
rect 11609 28948 11621 28951
rect 11480 28920 11621 28948
rect 11480 28908 11486 28920
rect 11609 28917 11621 28920
rect 11655 28917 11667 28951
rect 11609 28911 11667 28917
rect 17034 28908 17040 28960
rect 17092 28948 17098 28960
rect 19444 28948 19472 28988
rect 19886 28976 19892 28988
rect 19944 28976 19950 29028
rect 23293 29019 23351 29025
rect 23293 28985 23305 29019
rect 23339 29016 23351 29019
rect 23842 29016 23848 29028
rect 23339 28988 23848 29016
rect 23339 28985 23351 28988
rect 23293 28979 23351 28985
rect 23842 28976 23848 28988
rect 23900 29016 23906 29028
rect 24489 29019 24547 29025
rect 24489 29016 24501 29019
rect 23900 28988 24501 29016
rect 23900 28976 23906 28988
rect 24489 28985 24501 28988
rect 24535 28985 24547 29019
rect 24489 28979 24547 28985
rect 17092 28920 19472 28948
rect 17092 28908 17098 28920
rect 19518 28908 19524 28960
rect 19576 28948 19582 28960
rect 19797 28951 19855 28957
rect 19797 28948 19809 28951
rect 19576 28920 19809 28948
rect 19576 28908 19582 28920
rect 19797 28917 19809 28920
rect 19843 28917 19855 28951
rect 19797 28911 19855 28917
rect 24026 28908 24032 28960
rect 24084 28908 24090 28960
rect 1104 28858 28888 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 28888 28858
rect 1104 28784 28888 28806
rect 8665 28747 8723 28753
rect 8665 28744 8677 28747
rect 6886 28716 8677 28744
rect 5905 28679 5963 28685
rect 5905 28645 5917 28679
rect 5951 28676 5963 28679
rect 6886 28676 6914 28716
rect 8665 28713 8677 28716
rect 8711 28744 8723 28747
rect 10134 28744 10140 28756
rect 8711 28716 10140 28744
rect 8711 28713 8723 28716
rect 8665 28707 8723 28713
rect 10134 28704 10140 28716
rect 10192 28704 10198 28756
rect 11241 28747 11299 28753
rect 11241 28713 11253 28747
rect 11287 28744 11299 28747
rect 11330 28744 11336 28756
rect 11287 28716 11336 28744
rect 11287 28713 11299 28716
rect 11241 28707 11299 28713
rect 11330 28704 11336 28716
rect 11388 28704 11394 28756
rect 11609 28747 11667 28753
rect 11609 28713 11621 28747
rect 11655 28744 11667 28747
rect 12986 28744 12992 28756
rect 11655 28716 12992 28744
rect 11655 28713 11667 28716
rect 11609 28707 11667 28713
rect 5951 28648 6914 28676
rect 5951 28645 5963 28648
rect 5905 28639 5963 28645
rect 6380 28617 6408 28648
rect 11054 28636 11060 28688
rect 11112 28676 11118 28688
rect 11624 28676 11652 28707
rect 12986 28704 12992 28716
rect 13044 28704 13050 28756
rect 15286 28704 15292 28756
rect 15344 28744 15350 28756
rect 15933 28747 15991 28753
rect 15933 28744 15945 28747
rect 15344 28716 15945 28744
rect 15344 28704 15350 28716
rect 15933 28713 15945 28716
rect 15979 28713 15991 28747
rect 15933 28707 15991 28713
rect 16850 28704 16856 28756
rect 16908 28744 16914 28756
rect 17494 28744 17500 28756
rect 16908 28716 17500 28744
rect 16908 28704 16914 28716
rect 17494 28704 17500 28716
rect 17552 28744 17558 28756
rect 17773 28747 17831 28753
rect 17773 28744 17785 28747
rect 17552 28716 17785 28744
rect 17552 28704 17558 28716
rect 17773 28713 17785 28716
rect 17819 28713 17831 28747
rect 17773 28707 17831 28713
rect 26050 28704 26056 28756
rect 26108 28704 26114 28756
rect 11112 28648 11652 28676
rect 11112 28636 11118 28648
rect 17678 28636 17684 28688
rect 17736 28636 17742 28688
rect 21177 28679 21235 28685
rect 21177 28676 21189 28679
rect 20364 28648 21189 28676
rect 6365 28611 6423 28617
rect 6365 28577 6377 28611
rect 6411 28577 6423 28611
rect 6365 28571 6423 28577
rect 7929 28611 7987 28617
rect 7929 28577 7941 28611
rect 7975 28608 7987 28611
rect 9398 28608 9404 28620
rect 7975 28580 9404 28608
rect 7975 28577 7987 28580
rect 7929 28571 7987 28577
rect 9398 28568 9404 28580
rect 9456 28568 9462 28620
rect 9766 28608 9772 28620
rect 9600 28580 9772 28608
rect 4525 28543 4583 28549
rect 4525 28509 4537 28543
rect 4571 28540 4583 28543
rect 7745 28543 7803 28549
rect 4571 28512 5764 28540
rect 4571 28509 4583 28512
rect 4525 28503 4583 28509
rect 4798 28481 4804 28484
rect 4792 28472 4804 28481
rect 4759 28444 4804 28472
rect 4792 28435 4804 28444
rect 4798 28432 4804 28435
rect 4856 28432 4862 28484
rect 5736 28472 5764 28512
rect 7745 28509 7757 28543
rect 7791 28509 7803 28543
rect 7745 28503 7803 28509
rect 7190 28472 7196 28484
rect 5736 28444 7196 28472
rect 7190 28432 7196 28444
rect 7248 28432 7254 28484
rect 7285 28475 7343 28481
rect 7285 28441 7297 28475
rect 7331 28472 7343 28475
rect 7760 28472 7788 28503
rect 8294 28500 8300 28552
rect 8352 28540 8358 28552
rect 8389 28543 8447 28549
rect 8389 28540 8401 28543
rect 8352 28512 8401 28540
rect 8352 28500 8358 28512
rect 8389 28509 8401 28512
rect 8435 28509 8447 28543
rect 8389 28503 8447 28509
rect 8481 28543 8539 28549
rect 8481 28509 8493 28543
rect 8527 28540 8539 28543
rect 9600 28540 9628 28580
rect 9766 28568 9772 28580
rect 9824 28568 9830 28620
rect 9858 28568 9864 28620
rect 9916 28568 9922 28620
rect 13078 28568 13084 28620
rect 13136 28608 13142 28620
rect 20364 28617 20392 28648
rect 21177 28645 21189 28648
rect 21223 28645 21235 28679
rect 21177 28639 21235 28645
rect 15197 28611 15255 28617
rect 15197 28608 15209 28611
rect 13136 28580 15209 28608
rect 13136 28568 13142 28580
rect 15197 28577 15209 28580
rect 15243 28577 15255 28611
rect 15197 28571 15255 28577
rect 17313 28611 17371 28617
rect 17313 28577 17325 28611
rect 17359 28608 17371 28611
rect 17589 28611 17647 28617
rect 17589 28608 17601 28611
rect 17359 28580 17601 28608
rect 17359 28577 17371 28580
rect 17313 28571 17371 28577
rect 17589 28577 17601 28580
rect 17635 28577 17647 28611
rect 17589 28571 17647 28577
rect 20349 28611 20407 28617
rect 20349 28577 20361 28611
rect 20395 28577 20407 28611
rect 20349 28571 20407 28577
rect 21542 28568 21548 28620
rect 21600 28608 21606 28620
rect 21637 28611 21695 28617
rect 21637 28608 21649 28611
rect 21600 28580 21649 28608
rect 21600 28568 21606 28580
rect 21637 28577 21649 28580
rect 21683 28577 21695 28611
rect 21637 28571 21695 28577
rect 21729 28611 21787 28617
rect 21729 28577 21741 28611
rect 21775 28608 21787 28611
rect 23842 28608 23848 28620
rect 21775 28580 23848 28608
rect 21775 28577 21787 28580
rect 21729 28571 21787 28577
rect 8527 28512 9628 28540
rect 10128 28543 10186 28549
rect 8527 28509 8539 28512
rect 8481 28503 8539 28509
rect 10128 28509 10140 28543
rect 10174 28509 10186 28543
rect 10128 28503 10186 28509
rect 12069 28543 12127 28549
rect 12069 28509 12081 28543
rect 12115 28540 12127 28543
rect 14090 28540 14096 28552
rect 12115 28512 14096 28540
rect 12115 28509 12127 28512
rect 12069 28503 12127 28509
rect 7331 28444 8524 28472
rect 7331 28441 7343 28444
rect 7285 28435 7343 28441
rect 8496 28416 8524 28444
rect 8662 28432 8668 28484
rect 8720 28472 8726 28484
rect 9033 28475 9091 28481
rect 9033 28472 9045 28475
rect 8720 28444 9045 28472
rect 8720 28432 8726 28444
rect 9033 28441 9045 28444
rect 9079 28441 9091 28475
rect 9033 28435 9091 28441
rect 9122 28432 9128 28484
rect 9180 28472 9186 28484
rect 9217 28475 9275 28481
rect 9217 28472 9229 28475
rect 9180 28444 9229 28472
rect 9180 28432 9186 28444
rect 9217 28441 9229 28444
rect 9263 28441 9275 28475
rect 9217 28435 9275 28441
rect 10042 28432 10048 28484
rect 10100 28472 10106 28484
rect 10152 28472 10180 28503
rect 14090 28500 14096 28512
rect 14148 28500 14154 28552
rect 14185 28543 14243 28549
rect 14185 28509 14197 28543
rect 14231 28509 14243 28543
rect 14185 28503 14243 28509
rect 14461 28543 14519 28549
rect 14461 28509 14473 28543
rect 14507 28509 14519 28543
rect 14461 28503 14519 28509
rect 12342 28481 12348 28484
rect 10100 28444 10180 28472
rect 10100 28432 10106 28444
rect 12336 28435 12348 28481
rect 12342 28432 12348 28435
rect 12400 28432 12406 28484
rect 13814 28432 13820 28484
rect 13872 28472 13878 28484
rect 14200 28472 14228 28503
rect 13872 28444 14228 28472
rect 13872 28432 13878 28444
rect 6822 28364 6828 28416
rect 6880 28404 6886 28416
rect 6917 28407 6975 28413
rect 6917 28404 6929 28407
rect 6880 28376 6929 28404
rect 6880 28364 6886 28376
rect 6917 28373 6929 28376
rect 6963 28373 6975 28407
rect 6917 28367 6975 28373
rect 7466 28364 7472 28416
rect 7524 28404 7530 28416
rect 7561 28407 7619 28413
rect 7561 28404 7573 28407
rect 7524 28376 7573 28404
rect 7524 28364 7530 28376
rect 7561 28373 7573 28376
rect 7607 28373 7619 28407
rect 7561 28367 7619 28373
rect 8202 28364 8208 28416
rect 8260 28364 8266 28416
rect 8478 28364 8484 28416
rect 8536 28364 8542 28416
rect 9306 28364 9312 28416
rect 9364 28364 9370 28416
rect 9398 28364 9404 28416
rect 9456 28364 9462 28416
rect 9585 28407 9643 28413
rect 9585 28373 9597 28407
rect 9631 28404 9643 28407
rect 9950 28404 9956 28416
rect 9631 28376 9956 28404
rect 9631 28373 9643 28376
rect 9585 28367 9643 28373
rect 9950 28364 9956 28376
rect 10008 28364 10014 28416
rect 13449 28407 13507 28413
rect 13449 28373 13461 28407
rect 13495 28404 13507 28407
rect 13630 28404 13636 28416
rect 13495 28376 13636 28404
rect 13495 28373 13507 28376
rect 13449 28367 13507 28373
rect 13630 28364 13636 28376
rect 13688 28404 13694 28416
rect 14476 28404 14504 28503
rect 14642 28500 14648 28552
rect 14700 28500 14706 28552
rect 16574 28500 16580 28552
rect 16632 28500 16638 28552
rect 16666 28500 16672 28552
rect 16724 28540 16730 28552
rect 16853 28543 16911 28549
rect 16853 28540 16865 28543
rect 16724 28512 16865 28540
rect 16724 28500 16730 28512
rect 16853 28509 16865 28512
rect 16899 28509 16911 28543
rect 16853 28503 16911 28509
rect 17126 28500 17132 28552
rect 17184 28500 17190 28552
rect 17770 28500 17776 28552
rect 17828 28540 17834 28552
rect 17865 28543 17923 28549
rect 17865 28540 17877 28543
rect 17828 28512 17877 28540
rect 17828 28500 17834 28512
rect 17865 28509 17877 28512
rect 17911 28509 17923 28543
rect 17865 28503 17923 28509
rect 19518 28500 19524 28552
rect 19576 28500 19582 28552
rect 19886 28500 19892 28552
rect 19944 28540 19950 28552
rect 21744 28540 21772 28571
rect 23842 28568 23848 28580
rect 23900 28568 23906 28620
rect 24854 28568 24860 28620
rect 24912 28608 24918 28620
rect 25409 28611 25467 28617
rect 25409 28608 25421 28611
rect 24912 28580 25421 28608
rect 24912 28568 24918 28580
rect 25409 28577 25421 28580
rect 25455 28577 25467 28611
rect 25409 28571 25467 28577
rect 19944 28512 21772 28540
rect 19944 28500 19950 28512
rect 23198 28500 23204 28552
rect 23256 28540 23262 28552
rect 23293 28543 23351 28549
rect 23293 28540 23305 28543
rect 23256 28512 23305 28540
rect 23256 28500 23262 28512
rect 23293 28509 23305 28512
rect 23339 28540 23351 28543
rect 23569 28543 23627 28549
rect 23569 28540 23581 28543
rect 23339 28512 23581 28540
rect 23339 28509 23351 28512
rect 23293 28503 23351 28509
rect 23569 28509 23581 28512
rect 23615 28540 23627 28543
rect 23658 28540 23664 28552
rect 23615 28512 23664 28540
rect 23615 28509 23627 28512
rect 23569 28503 23627 28509
rect 23658 28500 23664 28512
rect 23716 28500 23722 28552
rect 24486 28500 24492 28552
rect 24544 28540 24550 28552
rect 25041 28543 25099 28549
rect 25041 28540 25053 28543
rect 24544 28512 25053 28540
rect 24544 28500 24550 28512
rect 25041 28509 25053 28512
rect 25087 28509 25099 28543
rect 25041 28503 25099 28509
rect 14921 28475 14979 28481
rect 14921 28441 14933 28475
rect 14967 28472 14979 28475
rect 16945 28475 17003 28481
rect 16945 28472 16957 28475
rect 14967 28444 16957 28472
rect 14967 28441 14979 28444
rect 14921 28435 14979 28441
rect 16945 28441 16957 28444
rect 16991 28472 17003 28475
rect 17678 28472 17684 28484
rect 16991 28444 17684 28472
rect 16991 28441 17003 28444
rect 16945 28435 17003 28441
rect 17678 28432 17684 28444
rect 17736 28432 17742 28484
rect 23845 28475 23903 28481
rect 23845 28441 23857 28475
rect 23891 28472 23903 28475
rect 24578 28472 24584 28484
rect 23891 28444 24584 28472
rect 23891 28441 23903 28444
rect 23845 28435 23903 28441
rect 24578 28432 24584 28444
rect 24636 28432 24642 28484
rect 13688 28376 14504 28404
rect 13688 28364 13694 28376
rect 19426 28364 19432 28416
rect 19484 28364 19490 28416
rect 20898 28364 20904 28416
rect 20956 28364 20962 28416
rect 21542 28364 21548 28416
rect 21600 28364 21606 28416
rect 23474 28364 23480 28416
rect 23532 28404 23538 28416
rect 24489 28407 24547 28413
rect 24489 28404 24501 28407
rect 23532 28376 24501 28404
rect 23532 28364 23538 28376
rect 24489 28373 24501 28376
rect 24535 28373 24547 28407
rect 24489 28367 24547 28373
rect 1104 28314 28888 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 28888 28314
rect 1104 28240 28888 28262
rect 8478 28200 8484 28212
rect 6656 28172 8484 28200
rect 6656 28073 6684 28172
rect 8478 28160 8484 28172
rect 8536 28160 8542 28212
rect 10042 28160 10048 28212
rect 10100 28160 10106 28212
rect 10229 28203 10287 28209
rect 10229 28169 10241 28203
rect 10275 28200 10287 28203
rect 10502 28200 10508 28212
rect 10275 28172 10508 28200
rect 10275 28169 10287 28172
rect 10229 28163 10287 28169
rect 10502 28160 10508 28172
rect 10560 28160 10566 28212
rect 10870 28160 10876 28212
rect 10928 28160 10934 28212
rect 12989 28203 13047 28209
rect 12989 28169 13001 28203
rect 13035 28200 13047 28203
rect 13078 28200 13084 28212
rect 13035 28172 13084 28200
rect 13035 28169 13047 28172
rect 12989 28163 13047 28169
rect 13078 28160 13084 28172
rect 13136 28160 13142 28212
rect 15378 28160 15384 28212
rect 15436 28200 15442 28212
rect 16117 28203 16175 28209
rect 16117 28200 16129 28203
rect 15436 28172 16129 28200
rect 15436 28160 15442 28172
rect 16117 28169 16129 28172
rect 16163 28200 16175 28203
rect 16163 28172 16574 28200
rect 16163 28169 16175 28172
rect 16117 28163 16175 28169
rect 14093 28135 14151 28141
rect 14093 28132 14105 28135
rect 7116 28104 14105 28132
rect 6089 28067 6147 28073
rect 6089 28033 6101 28067
rect 6135 28064 6147 28067
rect 6641 28067 6699 28073
rect 6641 28064 6653 28067
rect 6135 28036 6653 28064
rect 6135 28033 6147 28036
rect 6089 28027 6147 28033
rect 6641 28033 6653 28036
rect 6687 28033 6699 28067
rect 6641 28027 6699 28033
rect 6822 28024 6828 28076
rect 6880 28024 6886 28076
rect 7116 27996 7144 28104
rect 14093 28101 14105 28104
rect 14139 28132 14151 28135
rect 14182 28132 14188 28144
rect 14139 28104 14188 28132
rect 14139 28101 14151 28104
rect 14093 28095 14151 28101
rect 14182 28092 14188 28104
rect 14240 28092 14246 28144
rect 7466 28073 7472 28076
rect 7460 28064 7472 28073
rect 7427 28036 7472 28064
rect 7460 28027 7472 28036
rect 7466 28024 7472 28027
rect 7524 28024 7530 28076
rect 9950 28024 9956 28076
rect 10008 28024 10014 28076
rect 10134 28024 10140 28076
rect 10192 28064 10198 28076
rect 10321 28067 10379 28073
rect 10321 28064 10333 28067
rect 10192 28036 10333 28064
rect 10192 28024 10198 28036
rect 10321 28033 10333 28036
rect 10367 28033 10379 28067
rect 10321 28027 10379 28033
rect 11054 28024 11060 28076
rect 11112 28024 11118 28076
rect 11609 28067 11667 28073
rect 11609 28064 11621 28067
rect 11164 28036 11621 28064
rect 6886 27968 7144 27996
rect 106 27888 112 27940
rect 164 27928 170 27940
rect 6886 27928 6914 27968
rect 7190 27956 7196 28008
rect 7248 27956 7254 28008
rect 9401 27999 9459 28005
rect 9401 27965 9413 27999
rect 9447 27965 9459 27999
rect 9401 27959 9459 27965
rect 10413 27999 10471 28005
rect 10413 27965 10425 27999
rect 10459 27965 10471 27999
rect 10413 27959 10471 27965
rect 164 27900 6914 27928
rect 8573 27931 8631 27937
rect 164 27888 170 27900
rect 8573 27897 8585 27931
rect 8619 27928 8631 27931
rect 8662 27928 8668 27940
rect 8619 27900 8668 27928
rect 8619 27897 8631 27900
rect 8573 27891 8631 27897
rect 8662 27888 8668 27900
rect 8720 27928 8726 27940
rect 9416 27928 9444 27959
rect 8720 27900 9444 27928
rect 10428 27928 10456 27959
rect 10962 27956 10968 28008
rect 11020 27996 11026 28008
rect 11164 27996 11192 28036
rect 11609 28033 11621 28036
rect 11655 28033 11667 28067
rect 11609 28027 11667 28033
rect 11876 28067 11934 28073
rect 11876 28033 11888 28067
rect 11922 28064 11934 28067
rect 12158 28064 12164 28076
rect 11922 28036 12164 28064
rect 11922 28033 11934 28036
rect 11876 28027 11934 28033
rect 12158 28024 12164 28036
rect 12216 28024 12222 28076
rect 12710 28024 12716 28076
rect 12768 28064 12774 28076
rect 13449 28067 13507 28073
rect 13449 28064 13461 28067
rect 12768 28036 13461 28064
rect 12768 28024 12774 28036
rect 13449 28033 13461 28036
rect 13495 28033 13507 28067
rect 13449 28027 13507 28033
rect 11020 27968 11192 27996
rect 11241 27999 11299 28005
rect 11020 27956 11026 27968
rect 11241 27965 11253 27999
rect 11287 27996 11299 27999
rect 11422 27996 11428 28008
rect 11287 27968 11428 27996
rect 11287 27965 11299 27968
rect 11241 27959 11299 27965
rect 11422 27956 11428 27968
rect 11480 27956 11486 28008
rect 13354 27956 13360 28008
rect 13412 27956 13418 28008
rect 10502 27928 10508 27940
rect 10428 27900 10508 27928
rect 8720 27888 8726 27900
rect 10502 27888 10508 27900
rect 10560 27928 10566 27940
rect 13817 27931 13875 27937
rect 10560 27900 11008 27928
rect 10560 27888 10566 27900
rect 6457 27863 6515 27869
rect 6457 27829 6469 27863
rect 6503 27860 6515 27863
rect 6730 27860 6736 27872
rect 6503 27832 6736 27860
rect 6503 27829 6515 27832
rect 6457 27823 6515 27829
rect 6730 27820 6736 27832
rect 6788 27820 6794 27872
rect 8846 27820 8852 27872
rect 8904 27820 8910 27872
rect 10597 27863 10655 27869
rect 10597 27829 10609 27863
rect 10643 27860 10655 27863
rect 10870 27860 10876 27872
rect 10643 27832 10876 27860
rect 10643 27829 10655 27832
rect 10597 27823 10655 27829
rect 10870 27820 10876 27832
rect 10928 27820 10934 27872
rect 10980 27860 11008 27900
rect 13817 27897 13829 27931
rect 13863 27928 13875 27931
rect 13998 27928 14004 27940
rect 13863 27900 14004 27928
rect 13863 27897 13875 27900
rect 13817 27891 13875 27897
rect 13998 27888 14004 27900
rect 14056 27888 14062 27940
rect 16546 27928 16574 28172
rect 16942 28160 16948 28212
rect 17000 28200 17006 28212
rect 17773 28203 17831 28209
rect 17773 28200 17785 28203
rect 17000 28172 17785 28200
rect 17000 28160 17006 28172
rect 17773 28169 17785 28172
rect 17819 28169 17831 28203
rect 22094 28200 22100 28212
rect 17773 28163 17831 28169
rect 22066 28160 22100 28200
rect 22152 28160 22158 28212
rect 24026 28160 24032 28212
rect 24084 28160 24090 28212
rect 24486 28160 24492 28212
rect 24544 28160 24550 28212
rect 24578 28160 24584 28212
rect 24636 28200 24642 28212
rect 25225 28203 25283 28209
rect 25225 28200 25237 28203
rect 24636 28172 25237 28200
rect 24636 28160 24642 28172
rect 25225 28169 25237 28172
rect 25271 28169 25283 28203
rect 25225 28163 25283 28169
rect 17144 28104 18000 28132
rect 16666 28024 16672 28076
rect 16724 28064 16730 28076
rect 17144 28073 17172 28104
rect 17972 28076 18000 28104
rect 16761 28067 16819 28073
rect 16761 28064 16773 28067
rect 16724 28036 16773 28064
rect 16724 28024 16730 28036
rect 16761 28033 16773 28036
rect 16807 28033 16819 28067
rect 16761 28027 16819 28033
rect 17129 28067 17187 28073
rect 17129 28033 17141 28067
rect 17175 28033 17187 28067
rect 17129 28027 17187 28033
rect 17497 28067 17555 28073
rect 17497 28033 17509 28067
rect 17543 28064 17555 28067
rect 17678 28064 17684 28076
rect 17543 28036 17684 28064
rect 17543 28033 17555 28036
rect 17497 28027 17555 28033
rect 17678 28024 17684 28036
rect 17736 28024 17742 28076
rect 17954 28024 17960 28076
rect 18012 28024 18018 28076
rect 20898 28024 20904 28076
rect 20956 28024 20962 28076
rect 21085 28067 21143 28073
rect 21085 28033 21097 28067
rect 21131 28033 21143 28067
rect 21085 28027 21143 28033
rect 21361 28067 21419 28073
rect 21361 28033 21373 28067
rect 21407 28064 21419 28067
rect 22066 28064 22094 28160
rect 24596 28132 24624 28160
rect 23308 28104 24624 28132
rect 21407 28036 22094 28064
rect 21407 28033 21419 28036
rect 21361 28027 21419 28033
rect 17402 27956 17408 28008
rect 17460 27996 17466 28008
rect 18141 27999 18199 28005
rect 18141 27996 18153 27999
rect 17460 27968 18153 27996
rect 17460 27956 17466 27968
rect 18141 27965 18153 27968
rect 18187 27965 18199 27999
rect 18141 27959 18199 27965
rect 20622 27956 20628 28008
rect 20680 27996 20686 28008
rect 21100 27996 21128 28027
rect 22186 28024 22192 28076
rect 22244 28064 22250 28076
rect 22741 28067 22799 28073
rect 22741 28064 22753 28067
rect 22244 28036 22753 28064
rect 22244 28024 22250 28036
rect 22741 28033 22753 28036
rect 22787 28064 22799 28067
rect 23106 28064 23112 28076
rect 22787 28036 23112 28064
rect 22787 28033 22799 28036
rect 22741 28027 22799 28033
rect 23106 28024 23112 28036
rect 23164 28024 23170 28076
rect 23308 28073 23336 28104
rect 23293 28067 23351 28073
rect 23293 28033 23305 28067
rect 23339 28033 23351 28067
rect 23293 28027 23351 28033
rect 23308 27996 23336 28027
rect 23474 28024 23480 28076
rect 23532 28024 23538 28076
rect 24026 28024 24032 28076
rect 24084 28064 24090 28076
rect 24121 28067 24179 28073
rect 24121 28064 24133 28067
rect 24084 28036 24133 28064
rect 24084 28024 24090 28036
rect 24121 28033 24133 28036
rect 24167 28064 24179 28067
rect 24857 28067 24915 28073
rect 24857 28064 24869 28067
rect 24167 28036 24869 28064
rect 24167 28033 24179 28036
rect 24121 28027 24179 28033
rect 24857 28033 24869 28036
rect 24903 28033 24915 28067
rect 24857 28027 24915 28033
rect 24946 28024 24952 28076
rect 25004 28024 25010 28076
rect 20680 27968 23336 27996
rect 20680 27956 20686 27968
rect 23842 27956 23848 28008
rect 23900 27956 23906 28008
rect 17218 27928 17224 27940
rect 16546 27900 17224 27928
rect 17218 27888 17224 27900
rect 17276 27888 17282 27940
rect 12342 27860 12348 27872
rect 10980 27832 12348 27860
rect 12342 27820 12348 27832
rect 12400 27820 12406 27872
rect 20898 27820 20904 27872
rect 20956 27820 20962 27872
rect 21453 27863 21511 27869
rect 21453 27829 21465 27863
rect 21499 27860 21511 27863
rect 21542 27860 21548 27872
rect 21499 27832 21548 27860
rect 21499 27829 21511 27832
rect 21453 27823 21511 27829
rect 21542 27820 21548 27832
rect 21600 27860 21606 27872
rect 22002 27860 22008 27872
rect 21600 27832 22008 27860
rect 21600 27820 21606 27832
rect 22002 27820 22008 27832
rect 22060 27820 22066 27872
rect 23474 27820 23480 27872
rect 23532 27820 23538 27872
rect 1104 27770 28888 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 28888 27770
rect 1104 27696 28888 27718
rect 8481 27659 8539 27665
rect 8481 27625 8493 27659
rect 8527 27656 8539 27659
rect 9306 27656 9312 27668
rect 8527 27628 9312 27656
rect 8527 27625 8539 27628
rect 8481 27619 8539 27625
rect 9306 27616 9312 27628
rect 9364 27656 9370 27668
rect 9401 27659 9459 27665
rect 9401 27656 9413 27659
rect 9364 27628 9413 27656
rect 9364 27616 9370 27628
rect 9401 27625 9413 27628
rect 9447 27625 9459 27659
rect 9401 27619 9459 27625
rect 12158 27616 12164 27668
rect 12216 27616 12222 27668
rect 12710 27616 12716 27668
rect 12768 27616 12774 27668
rect 14182 27616 14188 27668
rect 14240 27616 14246 27668
rect 17586 27656 17592 27668
rect 14844 27628 17592 27656
rect 7837 27591 7895 27597
rect 7837 27557 7849 27591
rect 7883 27588 7895 27591
rect 8294 27588 8300 27600
rect 7883 27560 8300 27588
rect 7883 27557 7895 27560
rect 7837 27551 7895 27557
rect 8294 27548 8300 27560
rect 8352 27548 8358 27600
rect 8665 27591 8723 27597
rect 8665 27557 8677 27591
rect 8711 27588 8723 27591
rect 8711 27560 10364 27588
rect 8711 27557 8723 27560
rect 8665 27551 8723 27557
rect 8386 27480 8392 27532
rect 8444 27520 8450 27532
rect 9398 27520 9404 27532
rect 8444 27492 9404 27520
rect 8444 27480 8450 27492
rect 9398 27480 9404 27492
rect 9456 27480 9462 27532
rect 10336 27529 10364 27560
rect 10321 27523 10379 27529
rect 10321 27489 10333 27523
rect 10367 27489 10379 27523
rect 10321 27483 10379 27489
rect 13078 27480 13084 27532
rect 13136 27520 13142 27532
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 13136 27492 13277 27520
rect 13136 27480 13142 27492
rect 13265 27489 13277 27492
rect 13311 27489 13323 27523
rect 13265 27483 13323 27489
rect 14090 27480 14096 27532
rect 14148 27520 14154 27532
rect 14844 27529 14872 27628
rect 17586 27616 17592 27628
rect 17644 27616 17650 27668
rect 17678 27616 17684 27668
rect 17736 27616 17742 27668
rect 22186 27616 22192 27668
rect 22244 27616 22250 27668
rect 24946 27616 24952 27668
rect 25004 27656 25010 27668
rect 25133 27659 25191 27665
rect 25133 27656 25145 27659
rect 25004 27628 25145 27656
rect 25004 27616 25010 27628
rect 25133 27625 25145 27628
rect 25179 27625 25191 27659
rect 25133 27619 25191 27625
rect 16485 27591 16543 27597
rect 16485 27557 16497 27591
rect 16531 27588 16543 27591
rect 16574 27588 16580 27600
rect 16531 27560 16580 27588
rect 16531 27557 16543 27560
rect 16485 27551 16543 27557
rect 16574 27548 16580 27560
rect 16632 27548 16638 27600
rect 17494 27548 17500 27600
rect 17552 27548 17558 27600
rect 24121 27591 24179 27597
rect 24121 27557 24133 27591
rect 24167 27588 24179 27591
rect 24167 27560 24532 27588
rect 24167 27557 24179 27560
rect 24121 27551 24179 27557
rect 14829 27523 14887 27529
rect 14829 27520 14841 27523
rect 14148 27492 14841 27520
rect 14148 27480 14154 27492
rect 14829 27489 14841 27492
rect 14875 27489 14887 27523
rect 14829 27483 14887 27489
rect 16758 27480 16764 27532
rect 16816 27520 16822 27532
rect 16945 27523 17003 27529
rect 16945 27520 16957 27523
rect 16816 27492 16957 27520
rect 16816 27480 16822 27492
rect 16945 27489 16957 27492
rect 16991 27489 17003 27523
rect 16945 27483 17003 27489
rect 17034 27480 17040 27532
rect 17092 27480 17098 27532
rect 24504 27529 24532 27560
rect 24489 27523 24547 27529
rect 24489 27489 24501 27523
rect 24535 27489 24547 27523
rect 24489 27483 24547 27489
rect 6457 27455 6515 27461
rect 6457 27421 6469 27455
rect 6503 27452 6515 27455
rect 7190 27452 7196 27464
rect 6503 27424 7196 27452
rect 6503 27421 6515 27424
rect 6457 27415 6515 27421
rect 7190 27412 7196 27424
rect 7248 27412 7254 27464
rect 8202 27412 8208 27464
rect 8260 27412 8266 27464
rect 8481 27455 8539 27461
rect 8481 27421 8493 27455
rect 8527 27452 8539 27455
rect 9122 27452 9128 27464
rect 8527 27424 9128 27452
rect 8527 27421 8539 27424
rect 8481 27415 8539 27421
rect 9122 27412 9128 27424
rect 9180 27412 9186 27464
rect 10042 27412 10048 27464
rect 10100 27412 10106 27464
rect 11054 27412 11060 27464
rect 11112 27452 11118 27464
rect 11517 27455 11575 27461
rect 11517 27452 11529 27455
rect 11112 27424 11529 27452
rect 11112 27412 11118 27424
rect 11517 27421 11529 27424
rect 11563 27421 11575 27455
rect 11517 27415 11575 27421
rect 16850 27412 16856 27464
rect 16908 27452 16914 27464
rect 17126 27452 17132 27464
rect 16908 27424 17132 27452
rect 16908 27412 16914 27424
rect 17126 27412 17132 27424
rect 17184 27452 17190 27464
rect 17184 27424 17908 27452
rect 17184 27412 17190 27424
rect 17880 27396 17908 27424
rect 18138 27412 18144 27464
rect 18196 27412 18202 27464
rect 20809 27455 20867 27461
rect 20809 27421 20821 27455
rect 20855 27452 20867 27455
rect 21450 27452 21456 27464
rect 20855 27424 21456 27452
rect 20855 27421 20867 27424
rect 20809 27415 20867 27421
rect 21450 27412 21456 27424
rect 21508 27452 21514 27464
rect 22741 27455 22799 27461
rect 22741 27452 22753 27455
rect 21508 27424 22753 27452
rect 21508 27412 21514 27424
rect 22741 27421 22753 27424
rect 22787 27421 22799 27455
rect 22741 27415 22799 27421
rect 23008 27455 23066 27461
rect 23008 27421 23020 27455
rect 23054 27452 23066 27455
rect 23474 27452 23480 27464
rect 23054 27424 23480 27452
rect 23054 27421 23066 27424
rect 23008 27415 23066 27421
rect 23474 27412 23480 27424
rect 23532 27412 23538 27464
rect 28442 27412 28448 27464
rect 28500 27412 28506 27464
rect 6730 27393 6736 27396
rect 6724 27384 6736 27393
rect 6691 27356 6736 27384
rect 6724 27347 6736 27356
rect 6730 27344 6736 27347
rect 6788 27344 6794 27396
rect 15096 27387 15154 27393
rect 15096 27353 15108 27387
rect 15142 27384 15154 27387
rect 15194 27384 15200 27396
rect 15142 27356 15200 27384
rect 15142 27353 15154 27356
rect 15096 27347 15154 27353
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 16224 27356 16574 27384
rect 10686 27276 10692 27328
rect 10744 27316 10750 27328
rect 16224 27325 16252 27356
rect 10965 27319 11023 27325
rect 10965 27316 10977 27319
rect 10744 27288 10977 27316
rect 10744 27276 10750 27288
rect 10965 27285 10977 27288
rect 11011 27285 11023 27319
rect 10965 27279 11023 27285
rect 16209 27319 16267 27325
rect 16209 27285 16221 27319
rect 16255 27285 16267 27319
rect 16546 27316 16574 27356
rect 16666 27344 16672 27396
rect 16724 27384 16730 27396
rect 17649 27387 17707 27393
rect 17649 27384 17661 27387
rect 16724 27356 17661 27384
rect 16724 27344 16730 27356
rect 17649 27353 17661 27356
rect 17695 27353 17707 27387
rect 17649 27347 17707 27353
rect 17862 27344 17868 27396
rect 17920 27344 17926 27396
rect 20898 27344 20904 27396
rect 20956 27384 20962 27396
rect 21054 27387 21112 27393
rect 21054 27384 21066 27387
rect 20956 27356 21066 27384
rect 20956 27344 20962 27356
rect 21054 27353 21066 27356
rect 21100 27353 21112 27387
rect 21054 27347 21112 27353
rect 16758 27316 16764 27328
rect 16546 27288 16764 27316
rect 16209 27279 16267 27285
rect 16758 27276 16764 27288
rect 16816 27276 16822 27328
rect 17126 27276 17132 27328
rect 17184 27316 17190 27328
rect 17770 27316 17776 27328
rect 17184 27288 17776 27316
rect 17184 27276 17190 27288
rect 17770 27276 17776 27288
rect 17828 27316 17834 27328
rect 18233 27319 18291 27325
rect 18233 27316 18245 27319
rect 17828 27288 18245 27316
rect 17828 27276 17834 27288
rect 18233 27285 18245 27288
rect 18279 27285 18291 27319
rect 18233 27279 18291 27285
rect 1104 27226 28888 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 28888 27226
rect 1104 27152 28888 27174
rect 8386 27072 8392 27124
rect 8444 27072 8450 27124
rect 10042 27072 10048 27124
rect 10100 27072 10106 27124
rect 11054 27072 11060 27124
rect 11112 27072 11118 27124
rect 12069 27115 12127 27121
rect 12069 27081 12081 27115
rect 12115 27112 12127 27115
rect 12342 27112 12348 27124
rect 12115 27084 12348 27112
rect 12115 27081 12127 27084
rect 12069 27075 12127 27081
rect 12342 27072 12348 27084
rect 12400 27072 12406 27124
rect 12805 27115 12863 27121
rect 12805 27081 12817 27115
rect 12851 27112 12863 27115
rect 12986 27112 12992 27124
rect 12851 27084 12992 27112
rect 12851 27081 12863 27084
rect 12805 27075 12863 27081
rect 7190 27044 7196 27056
rect 7024 27016 7196 27044
rect 7024 26985 7052 27016
rect 7190 27004 7196 27016
rect 7248 27044 7254 27056
rect 9858 27044 9864 27056
rect 7248 27016 9864 27044
rect 7248 27004 7254 27016
rect 7009 26979 7067 26985
rect 7009 26945 7021 26979
rect 7055 26945 7067 26979
rect 7009 26939 7067 26945
rect 7276 26979 7334 26985
rect 7276 26945 7288 26979
rect 7322 26976 7334 26979
rect 8110 26976 8116 26988
rect 7322 26948 8116 26976
rect 7322 26945 7334 26948
rect 7276 26939 7334 26945
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 8680 26985 8708 27016
rect 9858 27004 9864 27016
rect 9916 27004 9922 27056
rect 10686 27004 10692 27056
rect 10744 27004 10750 27056
rect 10781 27047 10839 27053
rect 10781 27013 10793 27047
rect 10827 27044 10839 27047
rect 11422 27044 11428 27056
rect 10827 27016 11428 27044
rect 10827 27013 10839 27016
rect 10781 27007 10839 27013
rect 11422 27004 11428 27016
rect 11480 27004 11486 27056
rect 12820 27044 12848 27075
rect 12986 27072 12992 27084
rect 13044 27072 13050 27124
rect 13449 27115 13507 27121
rect 13449 27081 13461 27115
rect 13495 27112 13507 27115
rect 16666 27112 16672 27124
rect 13495 27084 16672 27112
rect 13495 27081 13507 27084
rect 13449 27075 13507 27081
rect 16666 27072 16672 27084
rect 16724 27072 16730 27124
rect 17402 27072 17408 27124
rect 17460 27072 17466 27124
rect 22370 27072 22376 27124
rect 22428 27072 22434 27124
rect 24026 27112 24032 27124
rect 23124 27084 24032 27112
rect 13906 27044 13912 27056
rect 12268 27016 12848 27044
rect 13648 27016 13912 27044
rect 8938 26985 8944 26988
rect 8665 26979 8723 26985
rect 8665 26945 8677 26979
rect 8711 26945 8723 26979
rect 8665 26939 8723 26945
rect 8932 26939 8944 26985
rect 8938 26936 8944 26939
rect 8996 26936 9002 26988
rect 10502 26936 10508 26988
rect 10560 26936 10566 26988
rect 10870 26936 10876 26988
rect 10928 26936 10934 26988
rect 12268 26985 12296 27016
rect 12253 26979 12311 26985
rect 12253 26945 12265 26979
rect 12299 26945 12311 26979
rect 12253 26939 12311 26945
rect 12437 26979 12495 26985
rect 12437 26945 12449 26979
rect 12483 26976 12495 26979
rect 12710 26976 12716 26988
rect 12483 26948 12716 26976
rect 12483 26945 12495 26948
rect 12437 26939 12495 26945
rect 12710 26936 12716 26948
rect 12768 26936 12774 26988
rect 13078 26936 13084 26988
rect 13136 26976 13142 26988
rect 13648 26985 13676 27016
rect 13906 27004 13912 27016
rect 13964 27044 13970 27056
rect 14642 27044 14648 27056
rect 13964 27016 14648 27044
rect 13964 27004 13970 27016
rect 14642 27004 14648 27016
rect 14700 27004 14706 27056
rect 17420 27044 17448 27072
rect 16546 27016 17448 27044
rect 13265 26979 13323 26985
rect 13265 26976 13277 26979
rect 13136 26948 13277 26976
rect 13136 26936 13142 26948
rect 13265 26945 13277 26948
rect 13311 26945 13323 26979
rect 13265 26939 13323 26945
rect 13633 26979 13691 26985
rect 13633 26945 13645 26979
rect 13679 26945 13691 26979
rect 13633 26939 13691 26945
rect 13814 26936 13820 26988
rect 13872 26936 13878 26988
rect 13998 26936 14004 26988
rect 14056 26976 14062 26988
rect 14185 26979 14243 26985
rect 14185 26976 14197 26979
rect 14056 26948 14197 26976
rect 14056 26936 14062 26948
rect 14185 26945 14197 26948
rect 14231 26945 14243 26979
rect 14185 26939 14243 26945
rect 14734 26936 14740 26988
rect 14792 26936 14798 26988
rect 16393 26979 16451 26985
rect 16393 26945 16405 26979
rect 16439 26976 16451 26979
rect 16546 26976 16574 27016
rect 20254 27004 20260 27056
rect 20312 27044 20318 27056
rect 22189 27047 22247 27053
rect 22189 27044 22201 27047
rect 20312 27016 22201 27044
rect 20312 27004 20318 27016
rect 22189 27013 22201 27016
rect 22235 27013 22247 27047
rect 22189 27007 22247 27013
rect 22281 27047 22339 27053
rect 22281 27013 22293 27047
rect 22327 27044 22339 27047
rect 22388 27044 22416 27072
rect 23124 27053 23152 27084
rect 24026 27072 24032 27084
rect 24084 27072 24090 27124
rect 25130 27072 25136 27124
rect 25188 27072 25194 27124
rect 22327 27016 22416 27044
rect 23109 27047 23167 27053
rect 22327 27013 22339 27016
rect 22281 27007 22339 27013
rect 23109 27013 23121 27047
rect 23155 27013 23167 27047
rect 23109 27007 23167 27013
rect 23216 27016 23980 27044
rect 16439 26948 16574 26976
rect 16439 26945 16451 26948
rect 16393 26939 16451 26945
rect 16758 26936 16764 26988
rect 16816 26936 16822 26988
rect 17954 26936 17960 26988
rect 18012 26976 18018 26988
rect 18325 26979 18383 26985
rect 18325 26976 18337 26979
rect 18012 26948 18337 26976
rect 18012 26936 18018 26948
rect 18325 26945 18337 26948
rect 18371 26945 18383 26979
rect 18325 26939 18383 26945
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26945 18475 26979
rect 18417 26939 18475 26945
rect 14366 26868 14372 26920
rect 14424 26908 14430 26920
rect 15013 26911 15071 26917
rect 15013 26908 15025 26911
rect 14424 26880 15025 26908
rect 14424 26868 14430 26880
rect 15013 26877 15025 26880
rect 15059 26877 15071 26911
rect 15013 26871 15071 26877
rect 16301 26911 16359 26917
rect 16301 26877 16313 26911
rect 16347 26908 16359 26911
rect 16850 26908 16856 26920
rect 16347 26880 16856 26908
rect 16347 26877 16359 26880
rect 16301 26871 16359 26877
rect 16850 26868 16856 26880
rect 16908 26868 16914 26920
rect 17678 26868 17684 26920
rect 17736 26908 17742 26920
rect 18432 26908 18460 26939
rect 18598 26936 18604 26988
rect 18656 26936 18662 26988
rect 20622 26936 20628 26988
rect 20680 26976 20686 26988
rect 21913 26979 21971 26985
rect 21913 26976 21925 26979
rect 20680 26948 21925 26976
rect 20680 26936 20686 26948
rect 21913 26945 21925 26948
rect 21959 26945 21971 26979
rect 21913 26939 21971 26945
rect 22002 26936 22008 26988
rect 22060 26976 22066 26988
rect 22378 26979 22436 26985
rect 22378 26976 22390 26979
rect 22060 26948 22105 26976
rect 22296 26948 22390 26976
rect 22060 26936 22066 26948
rect 22296 26920 22324 26948
rect 22378 26945 22390 26948
rect 22424 26945 22436 26979
rect 22833 26979 22891 26985
rect 22833 26976 22845 26979
rect 22378 26939 22436 26945
rect 22572 26948 22845 26976
rect 17736 26880 18460 26908
rect 17736 26868 17742 26880
rect 22278 26868 22284 26920
rect 22336 26868 22342 26920
rect 14461 26843 14519 26849
rect 14461 26809 14473 26843
rect 14507 26840 14519 26843
rect 17034 26840 17040 26852
rect 14507 26812 17040 26840
rect 14507 26809 14519 26812
rect 14461 26803 14519 26809
rect 17034 26800 17040 26812
rect 17092 26800 17098 26852
rect 22572 26849 22600 26948
rect 22833 26945 22845 26948
rect 22879 26945 22891 26979
rect 22833 26939 22891 26945
rect 23014 26936 23020 26988
rect 23072 26936 23078 26988
rect 23216 26985 23244 27016
rect 23952 26988 23980 27016
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26945 23259 26979
rect 23201 26939 23259 26945
rect 23753 26979 23811 26985
rect 23753 26945 23765 26979
rect 23799 26945 23811 26979
rect 23753 26939 23811 26945
rect 22557 26843 22615 26849
rect 22557 26809 22569 26843
rect 22603 26809 22615 26843
rect 22557 26803 22615 26809
rect 23385 26843 23443 26849
rect 23385 26809 23397 26843
rect 23431 26840 23443 26843
rect 23768 26840 23796 26939
rect 23934 26936 23940 26988
rect 23992 26936 23998 26988
rect 24026 26936 24032 26988
rect 24084 26936 24090 26988
rect 24305 26979 24363 26985
rect 24305 26945 24317 26979
rect 24351 26976 24363 26979
rect 25148 26976 25176 27072
rect 24351 26948 25176 26976
rect 24351 26945 24363 26948
rect 24305 26939 24363 26945
rect 25222 26936 25228 26988
rect 25280 26936 25286 26988
rect 24121 26911 24179 26917
rect 24121 26877 24133 26911
rect 24167 26877 24179 26911
rect 24121 26871 24179 26877
rect 24489 26911 24547 26917
rect 24489 26877 24501 26911
rect 24535 26908 24547 26911
rect 24857 26911 24915 26917
rect 24857 26908 24869 26911
rect 24535 26880 24869 26908
rect 24535 26877 24547 26880
rect 24489 26871 24547 26877
rect 24857 26877 24869 26880
rect 24903 26877 24915 26911
rect 24857 26871 24915 26877
rect 23431 26812 23796 26840
rect 24136 26840 24164 26871
rect 25222 26840 25228 26852
rect 24136 26812 25228 26840
rect 23431 26809 23443 26812
rect 23385 26803 23443 26809
rect 25222 26800 25228 26812
rect 25280 26800 25286 26852
rect 13630 26732 13636 26784
rect 13688 26732 13694 26784
rect 18785 26775 18843 26781
rect 18785 26741 18797 26775
rect 18831 26772 18843 26775
rect 19886 26772 19892 26784
rect 18831 26744 19892 26772
rect 18831 26741 18843 26744
rect 18785 26735 18843 26741
rect 19886 26732 19892 26744
rect 19944 26732 19950 26784
rect 24854 26732 24860 26784
rect 24912 26732 24918 26784
rect 24946 26732 24952 26784
rect 25004 26732 25010 26784
rect 1104 26682 28888 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 28888 26682
rect 1104 26608 28888 26630
rect 8110 26528 8116 26580
rect 8168 26528 8174 26580
rect 13814 26528 13820 26580
rect 13872 26528 13878 26580
rect 17678 26528 17684 26580
rect 17736 26528 17742 26580
rect 17954 26528 17960 26580
rect 18012 26528 18018 26580
rect 20622 26528 20628 26580
rect 20680 26528 20686 26580
rect 22649 26571 22707 26577
rect 22649 26537 22661 26571
rect 22695 26568 22707 26571
rect 23014 26568 23020 26580
rect 22695 26540 23020 26568
rect 22695 26537 22707 26540
rect 22649 26531 22707 26537
rect 23014 26528 23020 26540
rect 23072 26528 23078 26580
rect 8481 26435 8539 26441
rect 8481 26401 8493 26435
rect 8527 26432 8539 26435
rect 8846 26432 8852 26444
rect 8527 26404 8852 26432
rect 8527 26401 8539 26404
rect 8481 26395 8539 26401
rect 8846 26392 8852 26404
rect 8904 26392 8910 26444
rect 9398 26392 9404 26444
rect 9456 26432 9462 26444
rect 9585 26435 9643 26441
rect 9585 26432 9597 26435
rect 9456 26404 9597 26432
rect 9456 26392 9462 26404
rect 9585 26401 9597 26404
rect 9631 26401 9643 26435
rect 9585 26395 9643 26401
rect 18417 26435 18475 26441
rect 18417 26401 18429 26435
rect 18463 26432 18475 26435
rect 19150 26432 19156 26444
rect 18463 26404 19156 26432
rect 18463 26401 18475 26404
rect 18417 26395 18475 26401
rect 19150 26392 19156 26404
rect 19208 26392 19214 26444
rect 20162 26392 20168 26444
rect 20220 26392 20226 26444
rect 20254 26392 20260 26444
rect 20312 26392 20318 26444
rect 8294 26324 8300 26376
rect 8352 26324 8358 26376
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12437 26367 12495 26373
rect 12437 26364 12449 26367
rect 12308 26336 12449 26364
rect 12308 26324 12314 26336
rect 12437 26333 12449 26336
rect 12483 26333 12495 26367
rect 12437 26327 12495 26333
rect 17126 26324 17132 26376
rect 17184 26324 17190 26376
rect 17221 26367 17279 26373
rect 17221 26333 17233 26367
rect 17267 26333 17279 26367
rect 17221 26327 17279 26333
rect 17405 26367 17463 26373
rect 17405 26333 17417 26367
rect 17451 26333 17463 26367
rect 17405 26327 17463 26333
rect 17497 26367 17555 26373
rect 17497 26333 17509 26367
rect 17543 26364 17555 26367
rect 18138 26364 18144 26376
rect 17543 26336 18144 26364
rect 17543 26333 17555 26336
rect 17497 26327 17555 26333
rect 12710 26305 12716 26308
rect 12704 26259 12716 26305
rect 12710 26256 12716 26259
rect 12768 26256 12774 26308
rect 17034 26256 17040 26308
rect 17092 26296 17098 26308
rect 17236 26296 17264 26327
rect 17092 26268 17264 26296
rect 17420 26296 17448 26327
rect 18138 26324 18144 26336
rect 18196 26324 18202 26376
rect 18233 26367 18291 26373
rect 18233 26333 18245 26367
rect 18279 26333 18291 26367
rect 18233 26327 18291 26333
rect 18509 26367 18567 26373
rect 18509 26333 18521 26367
rect 18555 26364 18567 26367
rect 19426 26364 19432 26376
rect 18555 26336 19432 26364
rect 18555 26333 18567 26336
rect 18509 26327 18567 26333
rect 17862 26296 17868 26308
rect 17420 26268 17868 26296
rect 17092 26256 17098 26268
rect 17862 26256 17868 26268
rect 17920 26296 17926 26308
rect 18248 26296 18276 26327
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 19886 26324 19892 26376
rect 19944 26324 19950 26376
rect 20073 26367 20131 26373
rect 20073 26333 20085 26367
rect 20119 26333 20131 26367
rect 20073 26327 20131 26333
rect 20441 26367 20499 26373
rect 20441 26333 20453 26367
rect 20487 26364 20499 26367
rect 22002 26364 22008 26376
rect 20487 26336 22008 26364
rect 20487 26333 20499 26336
rect 20441 26327 20499 26333
rect 17920 26268 18276 26296
rect 20088 26296 20116 26327
rect 22002 26324 22008 26336
rect 22060 26324 22066 26376
rect 22370 26324 22376 26376
rect 22428 26364 22434 26376
rect 22465 26367 22523 26373
rect 22465 26364 22477 26367
rect 22428 26336 22477 26364
rect 22428 26324 22434 26336
rect 22465 26333 22477 26336
rect 22511 26333 22523 26367
rect 22465 26327 22523 26333
rect 21174 26296 21180 26308
rect 20088 26268 21180 26296
rect 17920 26256 17926 26268
rect 21174 26256 21180 26268
rect 21232 26256 21238 26308
rect 22278 26256 22284 26308
rect 22336 26296 22342 26308
rect 22830 26296 22836 26308
rect 22336 26268 22836 26296
rect 22336 26256 22342 26268
rect 22830 26256 22836 26268
rect 22888 26256 22894 26308
rect 9033 26231 9091 26237
rect 9033 26197 9045 26231
rect 9079 26228 9091 26231
rect 9306 26228 9312 26240
rect 9079 26200 9312 26228
rect 9079 26197 9091 26200
rect 9033 26191 9091 26197
rect 9306 26188 9312 26200
rect 9364 26188 9370 26240
rect 1104 26138 28888 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 28888 26138
rect 1104 26064 28888 26086
rect 8938 25984 8944 26036
rect 8996 26024 9002 26036
rect 9033 26027 9091 26033
rect 9033 26024 9045 26027
rect 8996 25996 9045 26024
rect 8996 25984 9002 25996
rect 9033 25993 9045 25996
rect 9079 25993 9091 26027
rect 9033 25987 9091 25993
rect 12710 25984 12716 26036
rect 12768 25984 12774 26036
rect 13354 26024 13360 26036
rect 13096 25996 13360 26024
rect 9217 25891 9275 25897
rect 9217 25857 9229 25891
rect 9263 25857 9275 25891
rect 9217 25851 9275 25857
rect 8294 25644 8300 25696
rect 8352 25684 8358 25696
rect 8665 25687 8723 25693
rect 8665 25684 8677 25687
rect 8352 25656 8677 25684
rect 8352 25644 8358 25656
rect 8665 25653 8677 25656
rect 8711 25684 8723 25687
rect 9232 25684 9260 25851
rect 9306 25848 9312 25900
rect 9364 25848 9370 25900
rect 13096 25897 13124 25996
rect 13354 25984 13360 25996
rect 13412 25984 13418 26036
rect 18598 25984 18604 26036
rect 18656 26024 18662 26036
rect 18785 26027 18843 26033
rect 18785 26024 18797 26027
rect 18656 25996 18797 26024
rect 18656 25984 18662 25996
rect 18785 25993 18797 25996
rect 18831 25993 18843 26027
rect 20990 26024 20996 26036
rect 18785 25987 18843 25993
rect 18984 25996 20996 26024
rect 18984 25897 19012 25996
rect 20990 25984 20996 25996
rect 21048 26024 21054 26036
rect 21174 26024 21180 26036
rect 21048 25996 21180 26024
rect 21048 25984 21054 25996
rect 21174 25984 21180 25996
rect 21232 25984 21238 26036
rect 19061 25959 19119 25965
rect 19061 25925 19073 25959
rect 19107 25956 19119 25959
rect 20162 25956 20168 25968
rect 19107 25928 20168 25956
rect 19107 25925 19119 25928
rect 19061 25919 19119 25925
rect 20162 25916 20168 25928
rect 20220 25916 20226 25968
rect 12897 25891 12955 25897
rect 12897 25888 12909 25891
rect 12452 25860 12909 25888
rect 9766 25684 9772 25696
rect 8711 25656 9772 25684
rect 8711 25653 8723 25656
rect 8665 25647 8723 25653
rect 9766 25644 9772 25656
rect 9824 25684 9830 25696
rect 12452 25693 12480 25860
rect 12897 25857 12909 25860
rect 12943 25857 12955 25891
rect 12897 25851 12955 25857
rect 13081 25891 13139 25897
rect 13081 25857 13093 25891
rect 13127 25857 13139 25891
rect 13081 25851 13139 25857
rect 18969 25891 19027 25897
rect 18969 25857 18981 25891
rect 19015 25857 19027 25891
rect 18969 25851 19027 25857
rect 19150 25848 19156 25900
rect 19208 25848 19214 25900
rect 19337 25891 19395 25897
rect 19337 25857 19349 25891
rect 19383 25888 19395 25891
rect 19426 25888 19432 25900
rect 19383 25860 19432 25888
rect 19383 25857 19395 25860
rect 19337 25851 19395 25857
rect 19426 25848 19432 25860
rect 19484 25848 19490 25900
rect 13906 25780 13912 25832
rect 13964 25780 13970 25832
rect 18598 25780 18604 25832
rect 18656 25820 18662 25832
rect 19168 25820 19196 25848
rect 18656 25792 19196 25820
rect 18656 25780 18662 25792
rect 25774 25780 25780 25832
rect 25832 25780 25838 25832
rect 12437 25687 12495 25693
rect 12437 25684 12449 25687
rect 9824 25656 12449 25684
rect 9824 25644 9830 25656
rect 12437 25653 12449 25656
rect 12483 25653 12495 25687
rect 12437 25647 12495 25653
rect 24946 25644 24952 25696
rect 25004 25684 25010 25696
rect 25222 25684 25228 25696
rect 25004 25656 25228 25684
rect 25004 25644 25010 25656
rect 25222 25644 25228 25656
rect 25280 25644 25286 25696
rect 1104 25594 28888 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 28888 25594
rect 1104 25520 28888 25542
rect 21085 25483 21143 25489
rect 21085 25449 21097 25483
rect 21131 25480 21143 25483
rect 21174 25480 21180 25492
rect 21131 25452 21180 25480
rect 21131 25449 21143 25452
rect 21085 25443 21143 25449
rect 21174 25440 21180 25452
rect 21232 25440 21238 25492
rect 19794 25236 19800 25288
rect 19852 25236 19858 25288
rect 19981 25279 20039 25285
rect 19981 25245 19993 25279
rect 20027 25276 20039 25279
rect 20530 25276 20536 25288
rect 20027 25248 20536 25276
rect 20027 25245 20039 25248
rect 19981 25239 20039 25245
rect 20530 25236 20536 25248
rect 20588 25236 20594 25288
rect 20898 25168 20904 25220
rect 20956 25168 20962 25220
rect 19518 25100 19524 25152
rect 19576 25140 19582 25152
rect 19889 25143 19947 25149
rect 19889 25140 19901 25143
rect 19576 25112 19901 25140
rect 19576 25100 19582 25112
rect 19889 25109 19901 25112
rect 19935 25109 19947 25143
rect 19889 25103 19947 25109
rect 20714 25100 20720 25152
rect 20772 25140 20778 25152
rect 21101 25143 21159 25149
rect 21101 25140 21113 25143
rect 20772 25112 21113 25140
rect 20772 25100 20778 25112
rect 21101 25109 21113 25112
rect 21147 25109 21159 25143
rect 21101 25103 21159 25109
rect 21266 25100 21272 25152
rect 21324 25100 21330 25152
rect 1104 25050 28888 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 28888 25050
rect 1104 24976 28888 24998
rect 18249 24939 18307 24945
rect 18249 24936 18261 24939
rect 18248 24905 18261 24936
rect 18295 24905 18307 24939
rect 18248 24899 18307 24905
rect 18046 24828 18052 24880
rect 18104 24828 18110 24880
rect 18248 24812 18276 24899
rect 21174 24868 21180 24880
rect 20364 24840 21180 24868
rect 12161 24803 12219 24809
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 12250 24800 12256 24812
rect 12207 24772 12256 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 12250 24760 12256 24772
rect 12308 24760 12314 24812
rect 12434 24809 12440 24812
rect 12428 24763 12440 24809
rect 12434 24760 12440 24763
rect 12492 24760 12498 24812
rect 18230 24760 18236 24812
rect 18288 24760 18294 24812
rect 19518 24760 19524 24812
rect 19576 24760 19582 24812
rect 20364 24800 20392 24840
rect 21174 24828 21180 24840
rect 21232 24868 21238 24880
rect 21545 24871 21603 24877
rect 21545 24868 21557 24871
rect 21232 24840 21557 24868
rect 21232 24828 21238 24840
rect 21545 24837 21557 24840
rect 21591 24837 21603 24871
rect 23382 24868 23388 24880
rect 21545 24831 21603 24837
rect 23124 24840 23388 24868
rect 20088 24772 20392 24800
rect 20441 24803 20499 24809
rect 20088 24744 20116 24772
rect 20441 24769 20453 24803
rect 20487 24800 20499 24803
rect 21082 24800 21088 24812
rect 20487 24772 21088 24800
rect 20487 24769 20499 24772
rect 20441 24763 20499 24769
rect 21082 24760 21088 24772
rect 21140 24760 21146 24812
rect 22094 24760 22100 24812
rect 22152 24760 22158 24812
rect 23124 24809 23152 24840
rect 23382 24828 23388 24840
rect 23440 24828 23446 24880
rect 23585 24871 23643 24877
rect 23585 24868 23597 24871
rect 23584 24837 23597 24868
rect 23631 24837 23643 24871
rect 23584 24831 23643 24837
rect 22833 24803 22891 24809
rect 22833 24769 22845 24803
rect 22879 24769 22891 24803
rect 22833 24763 22891 24769
rect 23109 24803 23167 24809
rect 23109 24769 23121 24803
rect 23155 24769 23167 24803
rect 23584 24800 23612 24831
rect 23750 24800 23756 24812
rect 23584 24772 23756 24800
rect 23109 24763 23167 24769
rect 19797 24735 19855 24741
rect 19797 24701 19809 24735
rect 19843 24732 19855 24735
rect 20070 24732 20076 24744
rect 19843 24704 20076 24732
rect 19843 24701 19855 24704
rect 19797 24695 19855 24701
rect 20070 24692 20076 24704
rect 20128 24692 20134 24744
rect 20165 24735 20223 24741
rect 20165 24701 20177 24735
rect 20211 24732 20223 24735
rect 20806 24732 20812 24744
rect 20211 24704 20812 24732
rect 20211 24701 20223 24704
rect 20165 24695 20223 24701
rect 20806 24692 20812 24704
rect 20864 24692 20870 24744
rect 20990 24692 20996 24744
rect 21048 24692 21054 24744
rect 22373 24735 22431 24741
rect 22373 24701 22385 24735
rect 22419 24701 22431 24735
rect 22848 24732 22876 24763
rect 23750 24760 23756 24772
rect 23808 24760 23814 24812
rect 24118 24732 24124 24744
rect 22848 24704 24124 24732
rect 22373 24695 22431 24701
rect 13541 24667 13599 24673
rect 13541 24633 13553 24667
rect 13587 24664 13599 24667
rect 13906 24664 13912 24676
rect 13587 24636 13912 24664
rect 13587 24633 13599 24636
rect 13541 24627 13599 24633
rect 13906 24624 13912 24636
rect 13964 24624 13970 24676
rect 18417 24667 18475 24673
rect 18417 24633 18429 24667
rect 18463 24664 18475 24667
rect 18506 24664 18512 24676
rect 18463 24636 18512 24664
rect 18463 24633 18475 24636
rect 18417 24627 18475 24633
rect 18506 24624 18512 24636
rect 18564 24664 18570 24676
rect 19705 24667 19763 24673
rect 19705 24664 19717 24667
rect 18564 24636 19717 24664
rect 18564 24624 18570 24636
rect 19705 24633 19717 24636
rect 19751 24664 19763 24667
rect 20714 24664 20720 24676
rect 19751 24636 20720 24664
rect 19751 24633 19763 24636
rect 19705 24627 19763 24633
rect 20714 24624 20720 24636
rect 20772 24624 20778 24676
rect 21266 24624 21272 24676
rect 21324 24664 21330 24676
rect 22281 24667 22339 24673
rect 22281 24664 22293 24667
rect 21324 24636 22293 24664
rect 21324 24624 21330 24636
rect 22281 24633 22293 24636
rect 22327 24633 22339 24667
rect 22388 24664 22416 24695
rect 24118 24692 24124 24704
rect 24176 24692 24182 24744
rect 22388 24636 23612 24664
rect 22281 24627 22339 24633
rect 23584 24608 23612 24636
rect 17954 24556 17960 24608
rect 18012 24596 18018 24608
rect 18233 24599 18291 24605
rect 18233 24596 18245 24599
rect 18012 24568 18245 24596
rect 18012 24556 18018 24568
rect 18233 24565 18245 24568
rect 18279 24565 18291 24599
rect 18233 24559 18291 24565
rect 19337 24599 19395 24605
rect 19337 24565 19349 24599
rect 19383 24596 19395 24599
rect 19426 24596 19432 24608
rect 19383 24568 19432 24596
rect 19383 24565 19395 24568
rect 19337 24559 19395 24565
rect 19426 24556 19432 24568
rect 19484 24556 19490 24608
rect 19794 24556 19800 24608
rect 19852 24596 19858 24608
rect 20257 24599 20315 24605
rect 20257 24596 20269 24599
rect 19852 24568 20269 24596
rect 19852 24556 19858 24568
rect 20257 24565 20269 24568
rect 20303 24565 20315 24599
rect 20257 24559 20315 24565
rect 20622 24556 20628 24608
rect 20680 24556 20686 24608
rect 21910 24556 21916 24608
rect 21968 24556 21974 24608
rect 22646 24556 22652 24608
rect 22704 24556 22710 24608
rect 23017 24599 23075 24605
rect 23017 24565 23029 24599
rect 23063 24596 23075 24599
rect 23106 24596 23112 24608
rect 23063 24568 23112 24596
rect 23063 24565 23075 24568
rect 23017 24559 23075 24565
rect 23106 24556 23112 24568
rect 23164 24556 23170 24608
rect 23566 24556 23572 24608
rect 23624 24556 23630 24608
rect 23753 24599 23811 24605
rect 23753 24565 23765 24599
rect 23799 24596 23811 24599
rect 24486 24596 24492 24608
rect 23799 24568 24492 24596
rect 23799 24565 23811 24568
rect 23753 24559 23811 24565
rect 24486 24556 24492 24568
rect 24544 24556 24550 24608
rect 1104 24506 28888 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 28888 24506
rect 1104 24432 28888 24454
rect 11977 24395 12035 24401
rect 11977 24361 11989 24395
rect 12023 24392 12035 24395
rect 12434 24392 12440 24404
rect 12023 24364 12440 24392
rect 12023 24361 12035 24364
rect 11977 24355 12035 24361
rect 12434 24352 12440 24364
rect 12492 24352 12498 24404
rect 20898 24352 20904 24404
rect 20956 24392 20962 24404
rect 21453 24395 21511 24401
rect 21453 24392 21465 24395
rect 20956 24364 21465 24392
rect 20956 24352 20962 24364
rect 21453 24361 21465 24364
rect 21499 24361 21511 24395
rect 21453 24355 21511 24361
rect 24670 24284 24676 24336
rect 24728 24324 24734 24336
rect 24765 24327 24823 24333
rect 24765 24324 24777 24327
rect 24728 24296 24777 24324
rect 24728 24284 24734 24296
rect 24765 24293 24777 24296
rect 24811 24293 24823 24327
rect 24765 24287 24823 24293
rect 17034 24216 17040 24268
rect 17092 24216 17098 24268
rect 18230 24256 18236 24268
rect 17696 24228 18236 24256
rect 842 24148 848 24200
rect 900 24188 906 24200
rect 1489 24191 1547 24197
rect 1489 24188 1501 24191
rect 900 24160 1501 24188
rect 900 24148 906 24160
rect 1489 24157 1501 24160
rect 1535 24157 1547 24191
rect 1489 24151 1547 24157
rect 11054 24148 11060 24200
rect 11112 24188 11118 24200
rect 11974 24188 11980 24200
rect 11112 24160 11980 24188
rect 11112 24148 11118 24160
rect 11974 24148 11980 24160
rect 12032 24148 12038 24200
rect 12618 24148 12624 24200
rect 12676 24148 12682 24200
rect 17494 24148 17500 24200
rect 17552 24148 17558 24200
rect 17586 24148 17592 24200
rect 17644 24188 17650 24200
rect 17696 24197 17724 24228
rect 18230 24216 18236 24228
rect 18288 24216 18294 24268
rect 20622 24216 20628 24268
rect 20680 24216 20686 24268
rect 22646 24216 22652 24268
rect 22704 24256 22710 24268
rect 23201 24259 23259 24265
rect 23201 24256 23213 24259
rect 22704 24228 23213 24256
rect 22704 24216 22710 24228
rect 23201 24225 23213 24228
rect 23247 24225 23259 24259
rect 23201 24219 23259 24225
rect 23566 24216 23572 24268
rect 23624 24256 23630 24268
rect 23937 24259 23995 24265
rect 23937 24256 23949 24259
rect 23624 24228 23949 24256
rect 23624 24216 23630 24228
rect 23937 24225 23949 24228
rect 23983 24225 23995 24259
rect 23937 24219 23995 24225
rect 17681 24191 17739 24197
rect 17681 24188 17693 24191
rect 17644 24160 17693 24188
rect 17644 24148 17650 24160
rect 17681 24157 17693 24160
rect 17727 24157 17739 24191
rect 17681 24151 17739 24157
rect 17773 24191 17831 24197
rect 17773 24157 17785 24191
rect 17819 24188 17831 24191
rect 18046 24188 18052 24200
rect 17819 24160 18052 24188
rect 17819 24157 17831 24160
rect 17773 24151 17831 24157
rect 17788 24120 17816 24151
rect 18046 24148 18052 24160
rect 18104 24148 18110 24200
rect 18138 24148 18144 24200
rect 18196 24188 18202 24200
rect 18785 24191 18843 24197
rect 18785 24188 18797 24191
rect 18196 24160 18797 24188
rect 18196 24148 18202 24160
rect 18785 24157 18797 24160
rect 18831 24157 18843 24191
rect 18785 24151 18843 24157
rect 19334 24148 19340 24200
rect 19392 24148 19398 24200
rect 20254 24148 20260 24200
rect 20312 24188 20318 24200
rect 22097 24191 22155 24197
rect 22097 24188 22109 24191
rect 20312 24160 22109 24188
rect 20312 24148 20318 24160
rect 22097 24157 22109 24160
rect 22143 24157 22155 24191
rect 22097 24151 22155 24157
rect 23750 24148 23756 24200
rect 23808 24148 23814 24200
rect 24486 24148 24492 24200
rect 24544 24148 24550 24200
rect 16546 24092 17816 24120
rect 10413 24055 10471 24061
rect 10413 24021 10425 24055
rect 10459 24052 10471 24055
rect 10594 24052 10600 24064
rect 10459 24024 10600 24052
rect 10459 24021 10471 24024
rect 10413 24015 10471 24021
rect 10594 24012 10600 24024
rect 10652 24012 10658 24064
rect 16298 24012 16304 24064
rect 16356 24052 16362 24064
rect 16393 24055 16451 24061
rect 16393 24052 16405 24055
rect 16356 24024 16405 24052
rect 16356 24012 16362 24024
rect 16393 24021 16405 24024
rect 16439 24052 16451 24055
rect 16546 24052 16574 24092
rect 21266 24080 21272 24132
rect 21324 24120 21330 24132
rect 23768 24120 23796 24148
rect 21324 24092 23796 24120
rect 21324 24080 21330 24092
rect 24302 24080 24308 24132
rect 24360 24120 24366 24132
rect 24765 24123 24823 24129
rect 24765 24120 24777 24123
rect 24360 24092 24777 24120
rect 24360 24080 24366 24092
rect 24765 24089 24777 24092
rect 24811 24120 24823 24123
rect 25041 24123 25099 24129
rect 25041 24120 25053 24123
rect 24811 24092 25053 24120
rect 24811 24089 24823 24092
rect 24765 24083 24823 24089
rect 25041 24089 25053 24092
rect 25087 24089 25099 24123
rect 25041 24083 25099 24089
rect 16439 24024 16574 24052
rect 16439 24021 16451 24024
rect 16393 24015 16451 24021
rect 17310 24012 17316 24064
rect 17368 24012 17374 24064
rect 19518 24012 19524 24064
rect 19576 24052 19582 24064
rect 19981 24055 20039 24061
rect 19981 24052 19993 24055
rect 19576 24024 19993 24052
rect 19576 24012 19582 24024
rect 19981 24021 19993 24024
rect 20027 24021 20039 24055
rect 19981 24015 20039 24021
rect 21174 24012 21180 24064
rect 21232 24012 21238 24064
rect 22646 24012 22652 24064
rect 22704 24012 22710 24064
rect 23106 24012 23112 24064
rect 23164 24052 23170 24064
rect 23569 24055 23627 24061
rect 23569 24052 23581 24055
rect 23164 24024 23581 24052
rect 23164 24012 23170 24024
rect 23569 24021 23581 24024
rect 23615 24021 23627 24055
rect 23569 24015 23627 24021
rect 24581 24055 24639 24061
rect 24581 24021 24593 24055
rect 24627 24052 24639 24055
rect 24946 24052 24952 24064
rect 24627 24024 24952 24052
rect 24627 24021 24639 24024
rect 24581 24015 24639 24021
rect 24946 24012 24952 24024
rect 25004 24012 25010 24064
rect 1104 23962 28888 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 28888 23962
rect 1104 23888 28888 23910
rect 10045 23851 10103 23857
rect 10045 23817 10057 23851
rect 10091 23848 10103 23851
rect 11054 23848 11060 23860
rect 10091 23820 11060 23848
rect 10091 23817 10103 23820
rect 10045 23811 10103 23817
rect 11054 23808 11060 23820
rect 11112 23808 11118 23860
rect 12066 23808 12072 23860
rect 12124 23848 12130 23860
rect 12253 23851 12311 23857
rect 12253 23848 12265 23851
rect 12124 23820 12265 23848
rect 12124 23808 12130 23820
rect 12253 23817 12265 23820
rect 12299 23817 12311 23851
rect 12253 23811 12311 23817
rect 16215 23851 16273 23857
rect 16215 23817 16227 23851
rect 16261 23848 16273 23851
rect 17494 23848 17500 23860
rect 16261 23820 17500 23848
rect 16261 23817 16273 23820
rect 16215 23811 16273 23817
rect 17494 23808 17500 23820
rect 17552 23808 17558 23860
rect 18138 23808 18144 23860
rect 18196 23808 18202 23860
rect 20073 23851 20131 23857
rect 20073 23817 20085 23851
rect 20119 23848 20131 23851
rect 20254 23848 20260 23860
rect 20119 23820 20260 23848
rect 20119 23817 20131 23820
rect 20073 23811 20131 23817
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 23477 23851 23535 23857
rect 23477 23817 23489 23851
rect 23523 23848 23535 23851
rect 23566 23848 23572 23860
rect 23523 23820 23572 23848
rect 23523 23817 23535 23820
rect 23477 23811 23535 23817
rect 23566 23808 23572 23820
rect 23624 23808 23630 23860
rect 25225 23851 25283 23857
rect 25225 23817 25237 23851
rect 25271 23848 25283 23851
rect 25774 23848 25780 23860
rect 25271 23820 25780 23848
rect 25271 23817 25283 23820
rect 25225 23811 25283 23817
rect 25774 23808 25780 23820
rect 25832 23808 25838 23860
rect 16298 23780 16304 23792
rect 10888 23752 13492 23780
rect 8754 23672 8760 23724
rect 8812 23712 8818 23724
rect 8921 23715 8979 23721
rect 8921 23712 8933 23715
rect 8812 23684 8933 23712
rect 8812 23672 8818 23684
rect 8921 23681 8933 23684
rect 8967 23681 8979 23715
rect 8921 23675 8979 23681
rect 9766 23672 9772 23724
rect 9824 23712 9830 23724
rect 10505 23715 10563 23721
rect 10505 23712 10517 23715
rect 9824 23684 10517 23712
rect 9824 23672 9830 23684
rect 10505 23681 10517 23684
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 8478 23604 8484 23656
rect 8536 23644 8542 23656
rect 8665 23647 8723 23653
rect 8665 23644 8677 23647
rect 8536 23616 8677 23644
rect 8536 23604 8542 23616
rect 8665 23613 8677 23616
rect 8711 23613 8723 23647
rect 10520 23644 10548 23675
rect 10594 23672 10600 23724
rect 10652 23672 10658 23724
rect 10888 23644 10916 23752
rect 11974 23672 11980 23724
rect 12032 23712 12038 23724
rect 12437 23715 12495 23721
rect 12437 23712 12449 23715
rect 12032 23684 12449 23712
rect 12032 23672 12038 23684
rect 12437 23681 12449 23684
rect 12483 23681 12495 23715
rect 12437 23675 12495 23681
rect 12529 23715 12587 23721
rect 12529 23681 12541 23715
rect 12575 23712 12587 23715
rect 12710 23712 12716 23724
rect 12575 23684 12716 23712
rect 12575 23681 12587 23684
rect 12529 23675 12587 23681
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 13464 23721 13492 23752
rect 15856 23752 16304 23780
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23712 13507 23715
rect 13909 23715 13967 23721
rect 13909 23712 13921 23715
rect 13495 23684 13921 23712
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 13909 23681 13921 23684
rect 13955 23712 13967 23715
rect 14458 23712 14464 23724
rect 13955 23684 14464 23712
rect 13955 23681 13967 23684
rect 13909 23675 13967 23681
rect 14458 23672 14464 23684
rect 14516 23672 14522 23724
rect 15657 23715 15715 23721
rect 15657 23681 15669 23715
rect 15703 23712 15715 23715
rect 15746 23712 15752 23724
rect 15703 23684 15752 23712
rect 15703 23681 15715 23684
rect 15657 23675 15715 23681
rect 15746 23672 15752 23684
rect 15804 23672 15810 23724
rect 15856 23721 15884 23752
rect 16298 23740 16304 23752
rect 16356 23740 16362 23792
rect 17028 23783 17086 23789
rect 17028 23749 17040 23783
rect 17074 23780 17086 23783
rect 17310 23780 17316 23792
rect 17074 23752 17316 23780
rect 17074 23749 17086 23752
rect 17028 23743 17086 23749
rect 17310 23740 17316 23752
rect 17368 23740 17374 23792
rect 19518 23740 19524 23792
rect 19576 23789 19582 23792
rect 19576 23780 19588 23789
rect 19576 23752 19621 23780
rect 19812 23752 21496 23780
rect 19576 23743 19588 23752
rect 19576 23740 19582 23743
rect 15841 23715 15899 23721
rect 15841 23681 15853 23715
rect 15887 23681 15899 23715
rect 15841 23675 15899 23681
rect 16117 23715 16175 23721
rect 16117 23681 16129 23715
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 16393 23715 16451 23721
rect 16393 23681 16405 23715
rect 16439 23712 16451 23715
rect 17586 23712 17592 23724
rect 16439 23684 17592 23712
rect 16439 23681 16451 23684
rect 16393 23675 16451 23681
rect 10520 23616 10916 23644
rect 8665 23607 8723 23613
rect 10888 23520 10916 23616
rect 12069 23647 12127 23653
rect 12069 23613 12081 23647
rect 12115 23613 12127 23647
rect 12069 23607 12127 23613
rect 12084 23576 12112 23607
rect 12158 23604 12164 23656
rect 12216 23604 12222 23656
rect 13265 23647 13323 23653
rect 13265 23613 13277 23647
rect 13311 23644 13323 23647
rect 14274 23644 14280 23656
rect 13311 23616 14280 23644
rect 13311 23613 13323 23616
rect 13265 23607 13323 23613
rect 14274 23604 14280 23616
rect 14332 23604 14338 23656
rect 15764 23644 15792 23672
rect 16132 23644 16160 23675
rect 17586 23672 17592 23684
rect 17644 23672 17650 23724
rect 19812 23721 19840 23752
rect 21468 23724 21496 23752
rect 19797 23715 19855 23721
rect 19797 23681 19809 23715
rect 19843 23681 19855 23715
rect 19797 23675 19855 23681
rect 21174 23672 21180 23724
rect 21232 23721 21238 23724
rect 21232 23712 21244 23721
rect 21232 23684 21277 23712
rect 21232 23675 21244 23684
rect 21232 23672 21238 23675
rect 21450 23672 21456 23724
rect 21508 23712 21514 23724
rect 23845 23715 23903 23721
rect 23845 23712 23857 23715
rect 21508 23684 23857 23712
rect 21508 23672 21514 23684
rect 23845 23681 23857 23684
rect 23891 23681 23903 23715
rect 23845 23675 23903 23681
rect 24112 23715 24170 23721
rect 24112 23681 24124 23715
rect 24158 23712 24170 23715
rect 24486 23712 24492 23724
rect 24158 23684 24492 23712
rect 24158 23681 24170 23684
rect 24112 23675 24170 23681
rect 24486 23672 24492 23684
rect 24544 23672 24550 23724
rect 15764 23616 16160 23644
rect 16758 23604 16764 23656
rect 16816 23604 16822 23656
rect 21910 23604 21916 23656
rect 21968 23644 21974 23656
rect 22465 23647 22523 23653
rect 22465 23644 22477 23647
rect 21968 23616 22477 23644
rect 21968 23604 21974 23616
rect 22465 23613 22477 23616
rect 22511 23613 22523 23647
rect 22465 23607 22523 23613
rect 22830 23604 22836 23656
rect 22888 23604 22894 23656
rect 13538 23576 13544 23588
rect 12084 23548 13544 23576
rect 13538 23536 13544 23548
rect 13596 23536 13602 23588
rect 842 23468 848 23520
rect 900 23508 906 23520
rect 1489 23511 1547 23517
rect 1489 23508 1501 23511
rect 900 23480 1501 23508
rect 900 23468 906 23480
rect 1489 23477 1501 23480
rect 1535 23477 1547 23511
rect 1489 23471 1547 23477
rect 10318 23468 10324 23520
rect 10376 23468 10382 23520
rect 10870 23468 10876 23520
rect 10928 23508 10934 23520
rect 10965 23511 11023 23517
rect 10965 23508 10977 23511
rect 10928 23480 10977 23508
rect 10928 23468 10934 23480
rect 10965 23477 10977 23480
rect 11011 23477 11023 23511
rect 10965 23471 11023 23477
rect 12713 23511 12771 23517
rect 12713 23477 12725 23511
rect 12759 23508 12771 23511
rect 13262 23508 13268 23520
rect 12759 23480 13268 23508
rect 12759 23477 12771 23480
rect 12713 23471 12771 23477
rect 13262 23468 13268 23480
rect 13320 23468 13326 23520
rect 13630 23468 13636 23520
rect 13688 23468 13694 23520
rect 15654 23468 15660 23520
rect 15712 23468 15718 23520
rect 18417 23511 18475 23517
rect 18417 23477 18429 23511
rect 18463 23508 18475 23511
rect 18598 23508 18604 23520
rect 18463 23480 18604 23508
rect 18463 23477 18475 23480
rect 18417 23471 18475 23477
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 21726 23468 21732 23520
rect 21784 23508 21790 23520
rect 21913 23511 21971 23517
rect 21913 23508 21925 23511
rect 21784 23480 21925 23508
rect 21784 23468 21790 23480
rect 21913 23477 21925 23480
rect 21959 23477 21971 23511
rect 21913 23471 21971 23477
rect 1104 23418 28888 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 28888 23418
rect 1104 23344 28888 23366
rect 11977 23307 12035 23313
rect 8588 23276 10640 23304
rect 8478 23168 8484 23180
rect 6886 23140 8484 23168
rect 5629 23103 5687 23109
rect 5629 23069 5641 23103
rect 5675 23100 5687 23103
rect 6454 23100 6460 23112
rect 5675 23072 6460 23100
rect 5675 23069 5687 23072
rect 5629 23063 5687 23069
rect 6454 23060 6460 23072
rect 6512 23100 6518 23112
rect 6886 23100 6914 23140
rect 8478 23128 8484 23140
rect 8536 23128 8542 23180
rect 6512 23072 6914 23100
rect 7837 23103 7895 23109
rect 6512 23060 6518 23072
rect 7837 23069 7849 23103
rect 7883 23100 7895 23103
rect 8588 23100 8616 23276
rect 10612 23236 10640 23276
rect 11977 23273 11989 23307
rect 12023 23304 12035 23307
rect 12158 23304 12164 23316
rect 12023 23276 12164 23304
rect 12023 23273 12035 23276
rect 11977 23267 12035 23273
rect 12158 23264 12164 23276
rect 12216 23264 12222 23316
rect 12618 23264 12624 23316
rect 12676 23304 12682 23316
rect 13725 23307 13783 23313
rect 13725 23304 13737 23307
rect 12676 23276 13737 23304
rect 12676 23264 12682 23276
rect 13725 23273 13737 23276
rect 13771 23273 13783 23307
rect 16758 23304 16764 23316
rect 13725 23267 13783 23273
rect 15580 23276 16764 23304
rect 12066 23236 12072 23248
rect 10612 23208 12072 23236
rect 12066 23196 12072 23208
rect 12124 23196 12130 23248
rect 12437 23239 12495 23245
rect 12437 23236 12449 23239
rect 12176 23208 12449 23236
rect 7883 23072 8616 23100
rect 7883 23069 7895 23072
rect 7837 23063 7895 23069
rect 4614 22992 4620 23044
rect 4672 23032 4678 23044
rect 5874 23035 5932 23041
rect 5874 23032 5886 23035
rect 4672 23004 5886 23032
rect 4672 22992 4678 23004
rect 5874 23001 5886 23004
rect 5920 23001 5932 23035
rect 5874 22995 5932 23001
rect 7009 22967 7067 22973
rect 7009 22933 7021 22967
rect 7055 22964 7067 22967
rect 7852 22964 7880 23063
rect 9398 23060 9404 23112
rect 9456 23100 9462 23112
rect 10597 23103 10655 23109
rect 10597 23100 10609 23103
rect 9456 23072 10609 23100
rect 9456 23060 9462 23072
rect 10597 23069 10609 23072
rect 10643 23069 10655 23103
rect 10597 23063 10655 23069
rect 11425 23103 11483 23109
rect 11425 23069 11437 23103
rect 11471 23100 11483 23103
rect 11790 23100 11796 23112
rect 11471 23072 11796 23100
rect 11471 23069 11483 23072
rect 11425 23063 11483 23069
rect 11790 23060 11796 23072
rect 11848 23060 11854 23112
rect 12176 23044 12204 23208
rect 12437 23205 12449 23208
rect 12483 23205 12495 23239
rect 12437 23199 12495 23205
rect 12529 23239 12587 23245
rect 12529 23205 12541 23239
rect 12575 23236 12587 23239
rect 12802 23236 12808 23248
rect 12575 23208 12808 23236
rect 12575 23205 12587 23208
rect 12529 23199 12587 23205
rect 12802 23196 12808 23208
rect 12860 23196 12866 23248
rect 13538 23196 13544 23248
rect 13596 23236 13602 23248
rect 14277 23239 14335 23245
rect 14277 23236 14289 23239
rect 13596 23208 14289 23236
rect 13596 23196 13602 23208
rect 14277 23205 14289 23208
rect 14323 23205 14335 23239
rect 14277 23199 14335 23205
rect 13722 23168 13728 23180
rect 12268 23140 13728 23168
rect 12268 23109 12296 23140
rect 13722 23128 13728 23140
rect 13780 23128 13786 23180
rect 13998 23128 14004 23180
rect 14056 23168 14062 23180
rect 15580 23177 15608 23276
rect 16758 23264 16764 23276
rect 16816 23304 16822 23316
rect 20717 23307 20775 23313
rect 16816 23276 18736 23304
rect 16816 23264 16822 23276
rect 16945 23239 17003 23245
rect 16945 23205 16957 23239
rect 16991 23236 17003 23239
rect 17034 23236 17040 23248
rect 16991 23208 17040 23236
rect 16991 23205 17003 23208
rect 16945 23199 17003 23205
rect 17034 23196 17040 23208
rect 17092 23196 17098 23248
rect 17957 23239 18015 23245
rect 17957 23205 17969 23239
rect 18003 23236 18015 23239
rect 18003 23208 18276 23236
rect 18003 23205 18015 23208
rect 17957 23199 18015 23205
rect 18248 23177 18276 23208
rect 15565 23171 15623 23177
rect 15565 23168 15577 23171
rect 14056 23140 15577 23168
rect 14056 23128 14062 23140
rect 15565 23137 15577 23140
rect 15611 23137 15623 23171
rect 15565 23131 15623 23137
rect 18233 23171 18291 23177
rect 18233 23137 18245 23171
rect 18279 23137 18291 23171
rect 18233 23131 18291 23137
rect 18708 23112 18736 23276
rect 20717 23273 20729 23307
rect 20763 23304 20775 23307
rect 20990 23304 20996 23316
rect 20763 23276 20996 23304
rect 20763 23273 20775 23276
rect 20717 23267 20775 23273
rect 20990 23264 20996 23276
rect 21048 23264 21054 23316
rect 21082 23264 21088 23316
rect 21140 23304 21146 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 21140 23276 21189 23304
rect 21140 23264 21146 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 22830 23264 22836 23316
rect 22888 23264 22894 23316
rect 23382 23264 23388 23316
rect 23440 23304 23446 23316
rect 23477 23307 23535 23313
rect 23477 23304 23489 23307
rect 23440 23276 23489 23304
rect 23440 23264 23446 23276
rect 23477 23273 23489 23276
rect 23523 23273 23535 23307
rect 23477 23267 23535 23273
rect 24486 23264 24492 23316
rect 24544 23264 24550 23316
rect 24578 23264 24584 23316
rect 24636 23304 24642 23316
rect 24857 23307 24915 23313
rect 24857 23304 24869 23307
rect 24636 23276 24869 23304
rect 24636 23264 24642 23276
rect 24857 23273 24869 23276
rect 24903 23273 24915 23307
rect 24857 23267 24915 23273
rect 21450 23168 21456 23180
rect 20364 23140 21456 23168
rect 12253 23103 12311 23109
rect 12253 23069 12265 23103
rect 12299 23069 12311 23103
rect 12253 23063 12311 23069
rect 12618 23060 12624 23112
rect 12676 23060 12682 23112
rect 12710 23060 12716 23112
rect 12768 23060 12774 23112
rect 13262 23060 13268 23112
rect 13320 23060 13326 23112
rect 13541 23103 13599 23109
rect 13541 23069 13553 23103
rect 13587 23069 13599 23103
rect 13541 23063 13599 23069
rect 10318 22992 10324 23044
rect 10376 23041 10382 23044
rect 10376 23032 10388 23041
rect 11701 23035 11759 23041
rect 10376 23004 10421 23032
rect 10376 22995 10388 23004
rect 11701 23001 11713 23035
rect 11747 23032 11759 23035
rect 12158 23032 12164 23044
rect 11747 23004 12164 23032
rect 11747 23001 11759 23004
rect 11701 22995 11759 23001
rect 10376 22992 10382 22995
rect 12158 22992 12164 23004
rect 12216 22992 12222 23044
rect 12989 23035 13047 23041
rect 12989 23001 13001 23035
rect 13035 23032 13047 23035
rect 13556 23032 13584 23063
rect 14458 23060 14464 23112
rect 14516 23060 14522 23112
rect 14642 23060 14648 23112
rect 14700 23060 14706 23112
rect 15654 23060 15660 23112
rect 15712 23100 15718 23112
rect 15821 23103 15879 23109
rect 15821 23100 15833 23103
rect 15712 23072 15833 23100
rect 15712 23060 15718 23072
rect 15821 23069 15833 23072
rect 15867 23069 15879 23103
rect 15821 23063 15879 23069
rect 17681 23103 17739 23109
rect 17681 23069 17693 23103
rect 17727 23100 17739 23103
rect 18138 23100 18144 23112
rect 17727 23072 18144 23100
rect 17727 23069 17739 23072
rect 17681 23063 17739 23069
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 18690 23060 18696 23112
rect 18748 23100 18754 23112
rect 19337 23103 19395 23109
rect 19337 23100 19349 23103
rect 18748 23072 19349 23100
rect 18748 23060 18754 23072
rect 19337 23069 19349 23072
rect 19383 23100 19395 23103
rect 20364 23100 20392 23140
rect 21450 23128 21456 23140
rect 21508 23128 21514 23180
rect 23934 23128 23940 23180
rect 23992 23168 23998 23180
rect 24029 23171 24087 23177
rect 24029 23168 24041 23171
rect 23992 23140 24041 23168
rect 23992 23128 23998 23140
rect 24029 23137 24041 23140
rect 24075 23137 24087 23171
rect 24029 23131 24087 23137
rect 24946 23128 24952 23180
rect 25004 23128 25010 23180
rect 19383 23072 20392 23100
rect 19383 23069 19395 23072
rect 19337 23063 19395 23069
rect 20530 23060 20536 23112
rect 20588 23100 20594 23112
rect 20993 23103 21051 23109
rect 20993 23100 21005 23103
rect 20588 23072 21005 23100
rect 20588 23060 20594 23072
rect 20993 23069 21005 23072
rect 21039 23069 21051 23103
rect 20993 23063 21051 23069
rect 21177 23103 21235 23109
rect 21177 23069 21189 23103
rect 21223 23100 21235 23103
rect 21266 23100 21272 23112
rect 21223 23072 21272 23100
rect 21223 23069 21235 23072
rect 21177 23063 21235 23069
rect 13035 23004 13584 23032
rect 14476 23032 14504 23060
rect 14921 23035 14979 23041
rect 14921 23032 14933 23035
rect 14476 23004 14933 23032
rect 13035 23001 13047 23004
rect 12989 22995 13047 23001
rect 14921 23001 14933 23004
rect 14967 23001 14979 23035
rect 14921 22995 14979 23001
rect 17954 22992 17960 23044
rect 18012 22992 18018 23044
rect 19426 22992 19432 23044
rect 19484 23032 19490 23044
rect 19582 23035 19640 23041
rect 19582 23032 19594 23035
rect 19484 23004 19594 23032
rect 19484 22992 19490 23004
rect 19582 23001 19594 23004
rect 19628 23001 19640 23035
rect 21008 23032 21036 23063
rect 21266 23060 21272 23072
rect 21324 23060 21330 23112
rect 21726 23109 21732 23112
rect 21720 23100 21732 23109
rect 21687 23072 21732 23100
rect 21720 23063 21732 23072
rect 21726 23060 21732 23063
rect 21784 23060 21790 23112
rect 24670 23060 24676 23112
rect 24728 23060 24734 23112
rect 23382 23032 23388 23044
rect 21008 23004 23388 23032
rect 19582 22995 19640 23001
rect 23382 22992 23388 23004
rect 23440 22992 23446 23044
rect 7055 22936 7880 22964
rect 7055 22933 7067 22936
rect 7009 22927 7067 22933
rect 8386 22924 8392 22976
rect 8444 22924 8450 22976
rect 9217 22967 9275 22973
rect 9217 22933 9229 22967
rect 9263 22964 9275 22967
rect 9766 22964 9772 22976
rect 9263 22936 9772 22964
rect 9263 22933 9275 22936
rect 9217 22927 9275 22933
rect 9766 22924 9772 22936
rect 9824 22964 9830 22976
rect 11606 22964 11612 22976
rect 9824 22936 11612 22964
rect 9824 22924 9830 22936
rect 11606 22924 11612 22936
rect 11664 22924 11670 22976
rect 11793 22967 11851 22973
rect 11793 22933 11805 22967
rect 11839 22964 11851 22967
rect 12342 22964 12348 22976
rect 11839 22936 12348 22964
rect 11839 22933 11851 22936
rect 11793 22927 11851 22933
rect 12342 22924 12348 22936
rect 12400 22924 12406 22976
rect 12526 22924 12532 22976
rect 12584 22964 12590 22976
rect 13357 22967 13415 22973
rect 13357 22964 13369 22967
rect 12584 22936 13369 22964
rect 12584 22924 12590 22936
rect 13357 22933 13369 22936
rect 13403 22933 13415 22967
rect 13357 22927 13415 22933
rect 17773 22967 17831 22973
rect 17773 22933 17785 22967
rect 17819 22964 17831 22967
rect 18046 22964 18052 22976
rect 17819 22936 18052 22964
rect 17819 22933 17831 22936
rect 17773 22927 17831 22933
rect 18046 22924 18052 22936
rect 18104 22924 18110 22976
rect 18414 22924 18420 22976
rect 18472 22964 18478 22976
rect 18877 22967 18935 22973
rect 18877 22964 18889 22967
rect 18472 22936 18889 22964
rect 18472 22924 18478 22936
rect 18877 22933 18889 22936
rect 18923 22933 18935 22967
rect 18877 22927 18935 22933
rect 1104 22874 28888 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 28888 22874
rect 1104 22800 28888 22822
rect 4614 22720 4620 22772
rect 4672 22720 4678 22772
rect 8665 22763 8723 22769
rect 8665 22729 8677 22763
rect 8711 22760 8723 22763
rect 8754 22760 8760 22772
rect 8711 22732 8760 22760
rect 8711 22729 8723 22732
rect 8665 22723 8723 22729
rect 8754 22720 8760 22732
rect 8812 22720 8818 22772
rect 12158 22720 12164 22772
rect 12216 22760 12222 22772
rect 12621 22763 12679 22769
rect 12621 22760 12633 22763
rect 12216 22732 12633 22760
rect 12216 22720 12222 22732
rect 12621 22729 12633 22732
rect 12667 22729 12679 22763
rect 12621 22723 12679 22729
rect 14274 22720 14280 22772
rect 14332 22720 14338 22772
rect 18509 22763 18567 22769
rect 18509 22729 18521 22763
rect 18555 22760 18567 22763
rect 19334 22760 19340 22772
rect 18555 22732 19340 22760
rect 18555 22729 18567 22732
rect 18509 22723 18567 22729
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 19794 22720 19800 22772
rect 19852 22720 19858 22772
rect 23753 22763 23811 22769
rect 23753 22729 23765 22763
rect 23799 22760 23811 22763
rect 23934 22760 23940 22772
rect 23799 22732 23940 22760
rect 23799 22729 23811 22732
rect 23753 22723 23811 22729
rect 23934 22720 23940 22732
rect 23992 22720 23998 22772
rect 24118 22720 24124 22772
rect 24176 22720 24182 22772
rect 13630 22652 13636 22704
rect 13688 22692 13694 22704
rect 13734 22695 13792 22701
rect 13734 22692 13746 22695
rect 13688 22664 13746 22692
rect 13688 22652 13694 22664
rect 13734 22661 13746 22664
rect 13780 22661 13792 22695
rect 13734 22655 13792 22661
rect 17954 22652 17960 22704
rect 18012 22692 18018 22704
rect 22646 22701 22652 22704
rect 18877 22695 18935 22701
rect 18877 22692 18889 22695
rect 18012 22664 18889 22692
rect 18012 22652 18018 22664
rect 18877 22661 18889 22664
rect 18923 22661 18935 22695
rect 22640 22692 22652 22701
rect 22607 22664 22652 22692
rect 18877 22655 18935 22661
rect 22640 22655 22652 22664
rect 22646 22652 22652 22655
rect 22704 22652 22710 22704
rect 24578 22692 24584 22704
rect 24044 22664 24584 22692
rect 4433 22627 4491 22633
rect 4433 22593 4445 22627
rect 4479 22624 4491 22627
rect 4614 22624 4620 22636
rect 4479 22596 4620 22624
rect 4479 22593 4491 22596
rect 4433 22587 4491 22593
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 8386 22584 8392 22636
rect 8444 22584 8450 22636
rect 8481 22627 8539 22633
rect 8481 22593 8493 22627
rect 8527 22593 8539 22627
rect 8481 22587 8539 22593
rect 4249 22559 4307 22565
rect 4249 22525 4261 22559
rect 4295 22556 4307 22559
rect 4985 22559 5043 22565
rect 4985 22556 4997 22559
rect 4295 22528 4997 22556
rect 4295 22525 4307 22528
rect 4249 22519 4307 22525
rect 4985 22525 4997 22528
rect 5031 22556 5043 22559
rect 5626 22556 5632 22568
rect 5031 22528 5632 22556
rect 5031 22525 5043 22528
rect 4985 22519 5043 22525
rect 5626 22516 5632 22528
rect 5684 22556 5690 22568
rect 8496 22556 8524 22587
rect 8570 22584 8576 22636
rect 8628 22624 8634 22636
rect 9398 22624 9404 22636
rect 8628 22596 9404 22624
rect 8628 22584 8634 22596
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 9668 22627 9726 22633
rect 9668 22593 9680 22627
rect 9714 22624 9726 22627
rect 10686 22624 10692 22636
rect 9714 22596 10692 22624
rect 9714 22593 9726 22596
rect 9668 22587 9726 22593
rect 10686 22584 10692 22596
rect 10744 22584 10750 22636
rect 12434 22584 12440 22636
rect 12492 22624 12498 22636
rect 12802 22624 12808 22636
rect 12492 22596 12808 22624
rect 12492 22584 12498 22596
rect 12802 22584 12808 22596
rect 12860 22624 12866 22636
rect 14829 22627 14887 22633
rect 14829 22624 14841 22627
rect 12860 22596 14841 22624
rect 12860 22584 12866 22596
rect 14829 22593 14841 22596
rect 14875 22593 14887 22627
rect 14829 22587 14887 22593
rect 18414 22584 18420 22636
rect 18472 22584 18478 22636
rect 18506 22584 18512 22636
rect 18564 22584 18570 22636
rect 18598 22584 18604 22636
rect 18656 22624 18662 22636
rect 19429 22627 19487 22633
rect 19429 22624 19441 22627
rect 18656 22596 19441 22624
rect 18656 22584 18662 22596
rect 19429 22593 19441 22596
rect 19475 22593 19487 22627
rect 19429 22587 19487 22593
rect 19981 22627 20039 22633
rect 19981 22593 19993 22627
rect 20027 22593 20039 22627
rect 19981 22587 20039 22593
rect 11790 22556 11796 22568
rect 5684 22528 9076 22556
rect 5684 22516 5690 22528
rect 9048 22429 9076 22528
rect 10796 22528 11796 22556
rect 10796 22497 10824 22528
rect 11790 22516 11796 22528
rect 11848 22556 11854 22568
rect 12161 22559 12219 22565
rect 12161 22556 12173 22559
rect 11848 22528 12173 22556
rect 11848 22516 11854 22528
rect 12161 22525 12173 22528
rect 12207 22525 12219 22559
rect 12161 22519 12219 22525
rect 13998 22516 14004 22568
rect 14056 22516 14062 22568
rect 18233 22559 18291 22565
rect 18233 22525 18245 22559
rect 18279 22525 18291 22559
rect 18524 22556 18552 22584
rect 19996 22556 20024 22587
rect 20070 22584 20076 22636
rect 20128 22584 20134 22636
rect 21450 22584 21456 22636
rect 21508 22624 21514 22636
rect 24044 22633 24072 22664
rect 24578 22652 24584 22664
rect 24636 22652 24642 22704
rect 22373 22627 22431 22633
rect 22373 22624 22385 22627
rect 21508 22596 22385 22624
rect 21508 22584 21514 22596
rect 22373 22593 22385 22596
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 24029 22627 24087 22633
rect 24029 22593 24041 22627
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22624 24271 22627
rect 24854 22624 24860 22636
rect 24259 22596 24860 22624
rect 24259 22593 24271 22596
rect 24213 22587 24271 22593
rect 18524 22528 20024 22556
rect 18233 22519 18291 22525
rect 10781 22491 10839 22497
rect 10781 22457 10793 22491
rect 10827 22457 10839 22491
rect 18248 22488 18276 22519
rect 23382 22516 23388 22568
rect 23440 22556 23446 22568
rect 24228 22556 24256 22587
rect 24854 22584 24860 22596
rect 24912 22584 24918 22636
rect 23440 22528 24256 22556
rect 23440 22516 23446 22528
rect 20530 22488 20536 22500
rect 18248 22460 20536 22488
rect 10781 22451 10839 22457
rect 20530 22448 20536 22460
rect 20588 22448 20594 22500
rect 9033 22423 9091 22429
rect 9033 22389 9045 22423
rect 9079 22420 9091 22423
rect 10870 22420 10876 22432
rect 9079 22392 10876 22420
rect 9079 22389 9091 22392
rect 9033 22383 9091 22389
rect 10870 22380 10876 22392
rect 10928 22420 10934 22432
rect 11149 22423 11207 22429
rect 11149 22420 11161 22423
rect 10928 22392 11161 22420
rect 10928 22380 10934 22392
rect 11149 22389 11161 22392
rect 11195 22389 11207 22423
rect 11149 22383 11207 22389
rect 11238 22380 11244 22432
rect 11296 22420 11302 22432
rect 11609 22423 11667 22429
rect 11609 22420 11621 22423
rect 11296 22392 11621 22420
rect 11296 22380 11302 22392
rect 11609 22389 11621 22392
rect 11655 22389 11667 22423
rect 11609 22383 11667 22389
rect 1104 22330 28888 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 28888 22330
rect 1104 22256 28888 22278
rect 10686 22176 10692 22228
rect 10744 22176 10750 22228
rect 12434 22176 12440 22228
rect 12492 22176 12498 22228
rect 14642 22176 14648 22228
rect 14700 22216 14706 22228
rect 14829 22219 14887 22225
rect 14829 22216 14841 22219
rect 14700 22188 14841 22216
rect 14700 22176 14706 22188
rect 14829 22185 14841 22188
rect 14875 22185 14887 22219
rect 14829 22179 14887 22185
rect 18690 22176 18696 22228
rect 18748 22176 18754 22228
rect 9766 22040 9772 22092
rect 9824 22040 9830 22092
rect 10413 22083 10471 22089
rect 10413 22049 10425 22083
rect 10459 22080 10471 22083
rect 11057 22083 11115 22089
rect 11057 22080 11069 22083
rect 10459 22052 11069 22080
rect 10459 22049 10471 22052
rect 10413 22043 10471 22049
rect 11057 22049 11069 22052
rect 11103 22049 11115 22083
rect 12526 22080 12532 22092
rect 11057 22043 11115 22049
rect 12084 22052 12532 22080
rect 1210 21972 1216 22024
rect 1268 22012 1274 22024
rect 1489 22015 1547 22021
rect 1489 22012 1501 22015
rect 1268 21984 1501 22012
rect 1268 21972 1274 21984
rect 1489 21981 1501 21984
rect 1535 22012 1547 22015
rect 1949 22015 2007 22021
rect 1949 22012 1961 22015
rect 1535 21984 1961 22012
rect 1535 21981 1547 21984
rect 1489 21975 1547 21981
rect 1949 21981 1961 21984
rect 1995 21981 2007 22015
rect 1949 21975 2007 21981
rect 10870 21972 10876 22024
rect 10928 21972 10934 22024
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 11882 22012 11888 22024
rect 11655 21984 11888 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 11882 21972 11888 21984
rect 11940 21972 11946 22024
rect 1673 21879 1731 21885
rect 1673 21845 1685 21879
rect 1719 21876 1731 21879
rect 4614 21876 4620 21888
rect 1719 21848 4620 21876
rect 1719 21845 1731 21848
rect 1673 21839 1731 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 12084 21876 12112 22052
rect 12526 22040 12532 22052
rect 12584 22040 12590 22092
rect 22094 22040 22100 22092
rect 22152 22080 22158 22092
rect 23201 22083 23259 22089
rect 23201 22080 23213 22083
rect 22152 22052 23213 22080
rect 22152 22040 22158 22052
rect 23201 22049 23213 22052
rect 23247 22049 23259 22083
rect 23201 22043 23259 22049
rect 12158 21972 12164 22024
rect 12216 22012 12222 22024
rect 13817 22015 13875 22021
rect 13817 22012 13829 22015
rect 12216 21984 13829 22012
rect 12216 21972 12222 21984
rect 13817 21981 13829 21984
rect 13863 22012 13875 22015
rect 13998 22012 14004 22024
rect 13863 21984 14004 22012
rect 13863 21981 13875 21984
rect 13817 21975 13875 21981
rect 13998 21972 14004 21984
rect 14056 21972 14062 22024
rect 14185 22015 14243 22021
rect 14185 21981 14197 22015
rect 14231 21981 14243 22015
rect 14185 21975 14243 21981
rect 13538 21904 13544 21956
rect 13596 21953 13602 21956
rect 13596 21907 13608 21953
rect 13596 21904 13602 21907
rect 13722 21904 13728 21956
rect 13780 21944 13786 21956
rect 14200 21944 14228 21975
rect 23106 21972 23112 22024
rect 23164 21972 23170 22024
rect 23293 22015 23351 22021
rect 23293 21981 23305 22015
rect 23339 22012 23351 22015
rect 23382 22012 23388 22024
rect 23339 21984 23388 22012
rect 23339 21981 23351 21984
rect 23293 21975 23351 21981
rect 23382 21972 23388 21984
rect 23440 21972 23446 22024
rect 17218 21944 17224 21956
rect 13780 21916 14228 21944
rect 16868 21916 17224 21944
rect 13780 21904 13786 21916
rect 16868 21888 16896 21916
rect 17218 21904 17224 21916
rect 17276 21904 17282 21956
rect 12161 21879 12219 21885
rect 12161 21876 12173 21879
rect 12084 21848 12173 21876
rect 12161 21845 12173 21848
rect 12207 21845 12219 21879
rect 12161 21839 12219 21845
rect 16850 21836 16856 21888
rect 16908 21836 16914 21888
rect 1104 21786 28888 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 28888 21786
rect 1104 21712 28888 21734
rect 12069 21675 12127 21681
rect 12069 21641 12081 21675
rect 12115 21672 12127 21675
rect 12618 21672 12624 21684
rect 12115 21644 12624 21672
rect 12115 21641 12127 21644
rect 12069 21635 12127 21641
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 11606 21564 11612 21616
rect 11664 21564 11670 21616
rect 10870 21496 10876 21548
rect 10928 21496 10934 21548
rect 11057 21539 11115 21545
rect 11057 21505 11069 21539
rect 11103 21536 11115 21539
rect 11238 21536 11244 21548
rect 11103 21508 11244 21536
rect 11103 21505 11115 21508
rect 11057 21499 11115 21505
rect 11238 21496 11244 21508
rect 11296 21496 11302 21548
rect 11790 21496 11796 21548
rect 11848 21496 11854 21548
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 11974 21536 11980 21548
rect 11931 21508 11980 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 12713 21539 12771 21545
rect 12713 21505 12725 21539
rect 12759 21536 12771 21539
rect 12894 21536 12900 21548
rect 12759 21508 12900 21536
rect 12759 21505 12771 21508
rect 12713 21499 12771 21505
rect 12894 21496 12900 21508
rect 12952 21536 12958 21548
rect 13446 21536 13452 21548
rect 12952 21508 13452 21536
rect 12952 21496 12958 21508
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 10413 21403 10471 21409
rect 10413 21369 10425 21403
rect 10459 21400 10471 21403
rect 10888 21400 10916 21496
rect 12250 21400 12256 21412
rect 10459 21372 12256 21400
rect 10459 21369 10471 21372
rect 10413 21363 10471 21369
rect 12250 21360 12256 21372
rect 12308 21400 12314 21412
rect 12308 21372 12434 21400
rect 12308 21360 12314 21372
rect 10689 21335 10747 21341
rect 10689 21301 10701 21335
rect 10735 21332 10747 21335
rect 10778 21332 10784 21344
rect 10735 21304 10784 21332
rect 10735 21301 10747 21304
rect 10689 21295 10747 21301
rect 10778 21292 10784 21304
rect 10836 21292 10842 21344
rect 11885 21335 11943 21341
rect 11885 21301 11897 21335
rect 11931 21332 11943 21335
rect 12066 21332 12072 21344
rect 11931 21304 12072 21332
rect 11931 21301 11943 21304
rect 11885 21295 11943 21301
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 12406 21332 12434 21372
rect 12621 21335 12679 21341
rect 12621 21332 12633 21335
rect 12406 21304 12633 21332
rect 12621 21301 12633 21304
rect 12667 21332 12679 21335
rect 13081 21335 13139 21341
rect 13081 21332 13093 21335
rect 12667 21304 13093 21332
rect 12667 21301 12679 21304
rect 12621 21295 12679 21301
rect 13081 21301 13093 21304
rect 13127 21301 13139 21335
rect 13081 21295 13139 21301
rect 1104 21242 28888 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 28888 21242
rect 1104 21168 28888 21190
rect 11882 21088 11888 21140
rect 11940 21088 11946 21140
rect 13541 21131 13599 21137
rect 13541 21097 13553 21131
rect 13587 21128 13599 21131
rect 13722 21128 13728 21140
rect 13587 21100 13728 21128
rect 13587 21097 13599 21100
rect 13541 21091 13599 21097
rect 13722 21088 13728 21100
rect 13780 21088 13786 21140
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 10505 20995 10563 21001
rect 10505 20992 10517 20995
rect 9456 20964 10517 20992
rect 9456 20952 9462 20964
rect 10505 20961 10517 20964
rect 10551 20961 10563 20995
rect 10505 20955 10563 20961
rect 12158 20952 12164 21004
rect 12216 20952 12222 21004
rect 15746 20992 15752 21004
rect 14936 20964 15752 20992
rect 10778 20933 10784 20936
rect 10772 20924 10784 20933
rect 10739 20896 10784 20924
rect 10772 20887 10784 20896
rect 10778 20884 10784 20887
rect 10836 20884 10842 20936
rect 14936 20933 14964 20964
rect 15746 20952 15752 20964
rect 15804 20952 15810 21004
rect 14921 20927 14979 20933
rect 14921 20893 14933 20927
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 15105 20927 15163 20933
rect 15105 20893 15117 20927
rect 15151 20893 15163 20927
rect 15105 20887 15163 20893
rect 12434 20865 12440 20868
rect 12428 20819 12440 20865
rect 12434 20816 12440 20819
rect 12492 20816 12498 20868
rect 15120 20856 15148 20887
rect 15562 20884 15568 20936
rect 15620 20884 15626 20936
rect 16209 20859 16267 20865
rect 16209 20856 16221 20859
rect 15120 20828 16221 20856
rect 16209 20825 16221 20828
rect 16255 20856 16267 20859
rect 16390 20856 16396 20868
rect 16255 20828 16396 20856
rect 16255 20825 16267 20828
rect 16209 20819 16267 20825
rect 16390 20816 16396 20828
rect 16448 20816 16454 20868
rect 15010 20748 15016 20800
rect 15068 20748 15074 20800
rect 1104 20698 28888 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 28888 20698
rect 1104 20624 28888 20646
rect 12434 20544 12440 20596
rect 12492 20544 12498 20596
rect 12526 20516 12532 20528
rect 12176 20488 12532 20516
rect 6454 20408 6460 20460
rect 6512 20408 6518 20460
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 12176 20457 12204 20488
rect 12526 20476 12532 20488
rect 12584 20476 12590 20528
rect 14820 20519 14878 20525
rect 14820 20485 14832 20519
rect 14866 20516 14878 20519
rect 15010 20516 15016 20528
rect 14866 20488 15016 20516
rect 14866 20485 14878 20488
rect 14820 20479 14878 20485
rect 15010 20476 15016 20488
rect 15068 20476 15074 20528
rect 19797 20519 19855 20525
rect 19797 20485 19809 20519
rect 19843 20485 19855 20519
rect 19797 20479 19855 20485
rect 6713 20451 6771 20457
rect 6713 20448 6725 20451
rect 6604 20420 6725 20448
rect 6604 20408 6610 20420
rect 6713 20417 6725 20420
rect 6759 20417 6771 20451
rect 6713 20411 6771 20417
rect 12161 20451 12219 20457
rect 12161 20417 12173 20451
rect 12207 20417 12219 20451
rect 12161 20411 12219 20417
rect 12250 20408 12256 20460
rect 12308 20448 12314 20460
rect 12713 20451 12771 20457
rect 12713 20448 12725 20451
rect 12308 20420 12725 20448
rect 12308 20408 12314 20420
rect 12713 20417 12725 20420
rect 12759 20417 12771 20451
rect 19812 20448 19840 20479
rect 19886 20476 19892 20528
rect 19944 20516 19950 20528
rect 19997 20519 20055 20525
rect 19997 20516 20009 20519
rect 19944 20488 20009 20516
rect 19944 20476 19950 20488
rect 19997 20485 20009 20488
rect 20043 20485 20055 20519
rect 19997 20479 20055 20485
rect 21818 20476 21824 20528
rect 21876 20516 21882 20528
rect 21913 20519 21971 20525
rect 21913 20516 21925 20519
rect 21876 20488 21925 20516
rect 21876 20476 21882 20488
rect 21913 20485 21925 20488
rect 21959 20485 21971 20519
rect 22113 20519 22171 20525
rect 22113 20516 22125 20519
rect 21913 20479 21971 20485
rect 22020 20488 22125 20516
rect 20254 20448 20260 20460
rect 19812 20420 20260 20448
rect 12713 20411 12771 20417
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 21174 20408 21180 20460
rect 21232 20448 21238 20460
rect 21269 20451 21327 20457
rect 21269 20448 21281 20451
rect 21232 20420 21281 20448
rect 21232 20408 21238 20420
rect 21269 20417 21281 20420
rect 21315 20448 21327 20451
rect 22020 20448 22048 20488
rect 22113 20485 22125 20488
rect 22159 20485 22171 20519
rect 22113 20479 22171 20485
rect 21315 20420 22048 20448
rect 22557 20451 22615 20457
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 22557 20417 22569 20451
rect 22603 20417 22615 20451
rect 22557 20411 22615 20417
rect 22741 20451 22799 20457
rect 22741 20417 22753 20451
rect 22787 20448 22799 20451
rect 22922 20448 22928 20460
rect 22787 20420 22928 20448
rect 22787 20417 22799 20420
rect 22741 20411 22799 20417
rect 13998 20340 14004 20392
rect 14056 20380 14062 20392
rect 14550 20380 14556 20392
rect 14056 20352 14556 20380
rect 14056 20340 14062 20352
rect 14550 20340 14556 20352
rect 14608 20340 14614 20392
rect 21082 20340 21088 20392
rect 21140 20340 21146 20392
rect 22572 20380 22600 20411
rect 22922 20408 22928 20420
rect 22980 20448 22986 20460
rect 23382 20448 23388 20460
rect 22980 20420 23388 20448
rect 22980 20408 22986 20420
rect 23382 20408 23388 20420
rect 23440 20408 23446 20460
rect 24486 20380 24492 20392
rect 22296 20352 24492 20380
rect 22002 20272 22008 20324
rect 22060 20312 22066 20324
rect 22296 20321 22324 20352
rect 24486 20340 24492 20352
rect 24544 20340 24550 20392
rect 22281 20315 22339 20321
rect 22060 20284 22140 20312
rect 22060 20272 22066 20284
rect 7837 20247 7895 20253
rect 7837 20213 7849 20247
rect 7883 20244 7895 20247
rect 8110 20244 8116 20256
rect 7883 20216 8116 20244
rect 7883 20213 7895 20216
rect 7837 20207 7895 20213
rect 8110 20204 8116 20216
rect 8168 20204 8174 20256
rect 15194 20204 15200 20256
rect 15252 20244 15258 20256
rect 15562 20244 15568 20256
rect 15252 20216 15568 20244
rect 15252 20204 15258 20216
rect 15562 20204 15568 20216
rect 15620 20244 15626 20256
rect 15933 20247 15991 20253
rect 15933 20244 15945 20247
rect 15620 20216 15945 20244
rect 15620 20204 15626 20216
rect 15933 20213 15945 20216
rect 15979 20213 15991 20247
rect 15933 20207 15991 20213
rect 19978 20204 19984 20256
rect 20036 20204 20042 20256
rect 20165 20247 20223 20253
rect 20165 20213 20177 20247
rect 20211 20244 20223 20247
rect 21174 20244 21180 20256
rect 20211 20216 21180 20244
rect 20211 20213 20223 20216
rect 20165 20207 20223 20213
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 21450 20204 21456 20256
rect 21508 20204 21514 20256
rect 22112 20253 22140 20284
rect 22281 20281 22293 20315
rect 22327 20281 22339 20315
rect 22281 20275 22339 20281
rect 22097 20247 22155 20253
rect 22097 20213 22109 20247
rect 22143 20213 22155 20247
rect 22097 20207 22155 20213
rect 22554 20204 22560 20256
rect 22612 20204 22618 20256
rect 1104 20154 28888 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 28888 20154
rect 1104 20080 28888 20102
rect 5626 20000 5632 20052
rect 5684 20000 5690 20052
rect 6365 20043 6423 20049
rect 6365 20009 6377 20043
rect 6411 20040 6423 20043
rect 6546 20040 6552 20052
rect 6411 20012 6552 20040
rect 6411 20009 6423 20012
rect 6365 20003 6423 20009
rect 6546 20000 6552 20012
rect 6604 20000 6610 20052
rect 18138 20000 18144 20052
rect 18196 20040 18202 20052
rect 18196 20012 18920 20040
rect 18196 20000 18202 20012
rect 5644 19904 5672 20000
rect 15562 19932 15568 19984
rect 15620 19972 15626 19984
rect 16209 19975 16267 19981
rect 16209 19972 16221 19975
rect 15620 19944 16221 19972
rect 15620 19932 15626 19944
rect 16209 19941 16221 19944
rect 16255 19941 16267 19975
rect 17773 19975 17831 19981
rect 17773 19972 17785 19975
rect 16209 19935 16267 19941
rect 16316 19944 17785 19972
rect 5644 19876 6224 19904
rect 6196 19845 6224 19876
rect 8110 19864 8116 19916
rect 8168 19864 8174 19916
rect 14550 19864 14556 19916
rect 14608 19864 14614 19916
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 16316 19904 16344 19944
rect 17773 19941 17785 19944
rect 17819 19972 17831 19975
rect 18892 19972 18920 20012
rect 21082 20000 21088 20052
rect 21140 20040 21146 20052
rect 22002 20040 22008 20052
rect 21140 20012 22008 20040
rect 21140 20000 21146 20012
rect 22002 20000 22008 20012
rect 22060 20040 22066 20052
rect 22465 20043 22523 20049
rect 22465 20040 22477 20043
rect 22060 20012 22477 20040
rect 22060 20000 22066 20012
rect 22465 20009 22477 20012
rect 22511 20009 22523 20043
rect 22465 20003 22523 20009
rect 23569 20043 23627 20049
rect 23569 20009 23581 20043
rect 23615 20040 23627 20043
rect 23658 20040 23664 20052
rect 23615 20012 23664 20040
rect 23615 20009 23627 20012
rect 23569 20003 23627 20009
rect 23658 20000 23664 20012
rect 23716 20040 23722 20052
rect 24302 20040 24308 20052
rect 23716 20012 24308 20040
rect 23716 20000 23722 20012
rect 24302 20000 24308 20012
rect 24360 20000 24366 20052
rect 21542 19972 21548 19984
rect 17819 19944 18828 19972
rect 18892 19944 21548 19972
rect 17819 19941 17831 19944
rect 17773 19935 17831 19941
rect 18233 19907 18291 19913
rect 18233 19904 18245 19907
rect 16080 19876 16344 19904
rect 17604 19876 18245 19904
rect 16080 19864 16086 19876
rect 6089 19839 6147 19845
rect 6089 19805 6101 19839
rect 6135 19805 6147 19839
rect 6089 19799 6147 19805
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19805 6239 19839
rect 6181 19799 6239 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 7834 19836 7840 19848
rect 7331 19808 7840 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 6104 19768 6132 19799
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 16390 19796 16396 19848
rect 16448 19796 16454 19848
rect 16482 19796 16488 19848
rect 16540 19796 16546 19848
rect 17604 19845 17632 19876
rect 18233 19873 18245 19876
rect 18279 19873 18291 19907
rect 18233 19867 18291 19873
rect 18800 19904 18828 19944
rect 21542 19932 21548 19944
rect 21600 19932 21606 19984
rect 19886 19904 19892 19916
rect 18800 19876 19892 19904
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19805 17647 19839
rect 17589 19799 17647 19805
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19805 17923 19839
rect 17865 19799 17923 19805
rect 6641 19771 6699 19777
rect 6641 19768 6653 19771
rect 6104 19740 6653 19768
rect 6641 19737 6653 19740
rect 6687 19768 6699 19771
rect 6730 19768 6736 19780
rect 6687 19740 6736 19768
rect 6687 19737 6699 19740
rect 6641 19731 6699 19737
rect 6730 19728 6736 19740
rect 6788 19728 6794 19780
rect 14820 19771 14878 19777
rect 14820 19737 14832 19771
rect 14866 19768 14878 19771
rect 15010 19768 15016 19780
rect 14866 19740 15016 19768
rect 14866 19737 14878 19740
rect 14820 19731 14878 19737
rect 15010 19728 15016 19740
rect 15068 19728 15074 19780
rect 15746 19728 15752 19780
rect 15804 19768 15810 19780
rect 16209 19771 16267 19777
rect 16209 19768 16221 19771
rect 15804 19740 16221 19768
rect 15804 19728 15810 19740
rect 16209 19737 16221 19740
rect 16255 19768 16267 19771
rect 17880 19768 17908 19799
rect 18138 19796 18144 19848
rect 18196 19796 18202 19848
rect 18322 19845 18328 19848
rect 18319 19799 18328 19845
rect 18380 19836 18386 19848
rect 18800 19845 18828 19876
rect 19886 19864 19892 19876
rect 19944 19864 19950 19916
rect 22922 19864 22928 19916
rect 22980 19864 22986 19916
rect 18785 19839 18843 19845
rect 18380 19808 18419 19836
rect 18322 19796 18328 19799
rect 18380 19796 18386 19808
rect 18785 19805 18797 19839
rect 18831 19805 18843 19839
rect 18785 19799 18843 19805
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 18892 19768 18920 19799
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 19521 19839 19579 19845
rect 19521 19836 19533 19839
rect 19024 19808 19533 19836
rect 19024 19796 19030 19808
rect 19521 19805 19533 19808
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 20809 19839 20867 19845
rect 20809 19805 20821 19839
rect 20855 19836 20867 19839
rect 21174 19836 21180 19848
rect 20855 19808 21180 19836
rect 20855 19805 20867 19808
rect 20809 19799 20867 19805
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21726 19796 21732 19848
rect 21784 19836 21790 19848
rect 21821 19839 21879 19845
rect 21821 19836 21833 19839
rect 21784 19808 21833 19836
rect 21784 19796 21790 19808
rect 21821 19805 21833 19808
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 22741 19839 22799 19845
rect 22741 19805 22753 19839
rect 22787 19836 22799 19839
rect 23658 19836 23664 19848
rect 22787 19808 23664 19836
rect 22787 19805 22799 19808
rect 22741 19799 22799 19805
rect 23658 19796 23664 19808
rect 23716 19796 23722 19848
rect 19978 19768 19984 19780
rect 16255 19740 17540 19768
rect 17880 19740 19984 19768
rect 16255 19737 16267 19740
rect 16209 19731 16267 19737
rect 7558 19660 7564 19712
rect 7616 19660 7622 19712
rect 15933 19703 15991 19709
rect 15933 19669 15945 19703
rect 15979 19700 15991 19703
rect 16298 19700 16304 19712
rect 15979 19672 16304 19700
rect 15979 19669 15991 19672
rect 15933 19663 15991 19669
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 17402 19660 17408 19712
rect 17460 19660 17466 19712
rect 17512 19700 17540 19740
rect 19978 19728 19984 19740
rect 20036 19768 20042 19780
rect 20165 19771 20223 19777
rect 20165 19768 20177 19771
rect 20036 19740 20177 19768
rect 20036 19728 20042 19740
rect 20165 19737 20177 19740
rect 20211 19737 20223 19771
rect 20165 19731 20223 19737
rect 18138 19700 18144 19712
rect 17512 19672 18144 19700
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 18322 19660 18328 19712
rect 18380 19700 18386 19712
rect 18601 19703 18659 19709
rect 18601 19700 18613 19703
rect 18380 19672 18613 19700
rect 18380 19660 18386 19672
rect 18601 19669 18613 19672
rect 18647 19700 18659 19703
rect 19426 19700 19432 19712
rect 18647 19672 19432 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 21358 19660 21364 19712
rect 21416 19660 21422 19712
rect 1104 19610 28888 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 28888 19610
rect 1104 19536 28888 19558
rect 7834 19456 7840 19508
rect 7892 19456 7898 19508
rect 13446 19456 13452 19508
rect 13504 19456 13510 19508
rect 15010 19456 15016 19508
rect 15068 19456 15074 19508
rect 19521 19499 19579 19505
rect 19521 19465 19533 19499
rect 19567 19496 19579 19499
rect 20898 19496 20904 19508
rect 19567 19468 20904 19496
rect 19567 19465 19579 19468
rect 19521 19459 19579 19465
rect 20898 19456 20904 19468
rect 20956 19496 20962 19508
rect 20956 19468 21312 19496
rect 20956 19456 20962 19468
rect 8972 19431 9030 19437
rect 8972 19397 8984 19431
rect 9018 19428 9030 19431
rect 10781 19431 10839 19437
rect 10781 19428 10793 19431
rect 9018 19400 10793 19428
rect 9018 19397 9030 19400
rect 8972 19391 9030 19397
rect 10781 19397 10793 19400
rect 10827 19428 10839 19431
rect 10870 19428 10876 19440
rect 10827 19400 10876 19428
rect 10827 19397 10839 19400
rect 10781 19391 10839 19397
rect 10870 19388 10876 19400
rect 10928 19388 10934 19440
rect 15746 19428 15752 19440
rect 13556 19400 15752 19428
rect 5629 19363 5687 19369
rect 5629 19360 5641 19363
rect 5460 19332 5641 19360
rect 4614 19252 4620 19304
rect 4672 19292 4678 19304
rect 5460 19292 5488 19332
rect 5629 19329 5641 19332
rect 5675 19360 5687 19363
rect 5902 19360 5908 19372
rect 5675 19332 5908 19360
rect 5675 19329 5687 19332
rect 5629 19323 5687 19329
rect 5902 19320 5908 19332
rect 5960 19320 5966 19372
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 9398 19360 9404 19372
rect 9263 19332 9404 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 10594 19320 10600 19372
rect 10652 19320 10658 19372
rect 13556 19369 13584 19400
rect 15746 19388 15752 19400
rect 15804 19388 15810 19440
rect 16390 19428 16396 19440
rect 15856 19400 16396 19428
rect 13541 19363 13599 19369
rect 13541 19329 13553 19363
rect 13587 19329 13599 19363
rect 13541 19323 13599 19329
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19360 15255 19363
rect 15562 19360 15568 19372
rect 15243 19332 15568 19360
rect 15243 19329 15255 19332
rect 15197 19323 15255 19329
rect 15562 19320 15568 19332
rect 15620 19320 15626 19372
rect 15856 19360 15884 19400
rect 16390 19388 16396 19400
rect 16448 19388 16454 19440
rect 15672 19332 15884 19360
rect 15672 19304 15700 19332
rect 16022 19320 16028 19372
rect 16080 19320 16086 19372
rect 16482 19360 16488 19372
rect 16224 19332 16488 19360
rect 16224 19304 16252 19332
rect 16482 19320 16488 19332
rect 16540 19360 16546 19372
rect 16761 19363 16819 19369
rect 16761 19360 16773 19363
rect 16540 19332 16773 19360
rect 16540 19320 16546 19332
rect 16761 19329 16773 19332
rect 16807 19329 16819 19363
rect 16761 19323 16819 19329
rect 18408 19363 18466 19369
rect 18408 19329 18420 19363
rect 18454 19360 18466 19363
rect 19797 19363 19855 19369
rect 19797 19360 19809 19363
rect 18454 19332 19809 19360
rect 18454 19329 18466 19332
rect 18408 19323 18466 19329
rect 19797 19329 19809 19332
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 20254 19320 20260 19372
rect 20312 19360 20318 19372
rect 21284 19369 21312 19468
rect 21818 19456 21824 19508
rect 21876 19496 21882 19508
rect 23293 19499 23351 19505
rect 23293 19496 23305 19499
rect 21876 19468 23305 19496
rect 21876 19456 21882 19468
rect 23293 19465 23305 19468
rect 23339 19465 23351 19499
rect 23293 19459 23351 19465
rect 24302 19456 24308 19508
rect 24360 19456 24366 19508
rect 21542 19388 21548 19440
rect 21600 19428 21606 19440
rect 21600 19400 22140 19428
rect 21600 19388 21606 19400
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20312 19332 20729 19360
rect 20312 19320 20318 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 21450 19320 21456 19372
rect 21508 19360 21514 19372
rect 21913 19363 21971 19369
rect 21913 19360 21925 19363
rect 21508 19332 21925 19360
rect 21508 19320 21514 19332
rect 21913 19329 21925 19332
rect 21959 19360 21971 19363
rect 22002 19360 22008 19372
rect 21959 19332 22008 19360
rect 21959 19329 21971 19332
rect 21913 19323 21971 19329
rect 22002 19320 22008 19332
rect 22060 19320 22066 19372
rect 22112 19369 22140 19400
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19360 22155 19363
rect 22922 19360 22928 19372
rect 22143 19332 22928 19360
rect 22143 19329 22155 19332
rect 22097 19323 22155 19329
rect 22922 19320 22928 19332
rect 22980 19320 22986 19372
rect 4672 19264 5488 19292
rect 5813 19295 5871 19301
rect 4672 19252 4678 19264
rect 5813 19261 5825 19295
rect 5859 19292 5871 19295
rect 6457 19295 6515 19301
rect 6457 19292 6469 19295
rect 5859 19264 6469 19292
rect 5859 19261 5871 19264
rect 5813 19255 5871 19261
rect 6457 19261 6469 19264
rect 6503 19261 6515 19295
rect 6457 19255 6515 19261
rect 7098 19252 7104 19304
rect 7156 19252 7162 19304
rect 10042 19252 10048 19304
rect 10100 19252 10106 19304
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19292 10471 19295
rect 10502 19292 10508 19304
rect 10459 19264 10508 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 10502 19252 10508 19264
rect 10560 19252 10566 19304
rect 15473 19295 15531 19301
rect 15473 19261 15485 19295
rect 15519 19292 15531 19295
rect 15654 19292 15660 19304
rect 15519 19264 15660 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 15654 19252 15660 19264
rect 15712 19252 15718 19304
rect 16206 19292 16212 19304
rect 15856 19264 16212 19292
rect 15381 19227 15439 19233
rect 15381 19193 15393 19227
rect 15427 19224 15439 19227
rect 15856 19224 15884 19264
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16298 19252 16304 19304
rect 16356 19292 16362 19304
rect 17313 19295 17371 19301
rect 17313 19292 17325 19295
rect 16356 19264 17325 19292
rect 16356 19252 16362 19264
rect 17313 19261 17325 19264
rect 17359 19261 17371 19295
rect 17313 19255 17371 19261
rect 18138 19252 18144 19304
rect 18196 19252 18202 19304
rect 20346 19252 20352 19304
rect 20404 19252 20410 19304
rect 22370 19252 22376 19304
rect 22428 19252 22434 19304
rect 23842 19252 23848 19304
rect 23900 19252 23906 19304
rect 15427 19196 15884 19224
rect 15933 19227 15991 19233
rect 15427 19193 15439 19196
rect 15381 19187 15439 19193
rect 15933 19193 15945 19227
rect 15979 19224 15991 19227
rect 16666 19224 16672 19236
rect 15979 19196 16672 19224
rect 15979 19193 15991 19196
rect 15933 19187 15991 19193
rect 16666 19184 16672 19196
rect 16724 19184 16730 19236
rect 5442 19116 5448 19168
rect 5500 19116 5506 19168
rect 9214 19116 9220 19168
rect 9272 19156 9278 19168
rect 9493 19159 9551 19165
rect 9493 19156 9505 19159
rect 9272 19128 9505 19156
rect 9272 19116 9278 19128
rect 9493 19125 9505 19128
rect 9539 19125 9551 19159
rect 9493 19119 9551 19125
rect 15838 19116 15844 19168
rect 15896 19116 15902 19168
rect 20990 19116 20996 19168
rect 21048 19156 21054 19168
rect 21913 19159 21971 19165
rect 21913 19156 21925 19159
rect 21048 19128 21925 19156
rect 21048 19116 21054 19128
rect 21913 19125 21925 19128
rect 21959 19125 21971 19159
rect 21913 19119 21971 19125
rect 23017 19159 23075 19165
rect 23017 19125 23029 19159
rect 23063 19156 23075 19159
rect 23106 19156 23112 19168
rect 23063 19128 23112 19156
rect 23063 19125 23075 19128
rect 23017 19119 23075 19125
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 1104 19066 28888 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 28888 19066
rect 1104 18992 28888 19014
rect 7098 18912 7104 18964
rect 7156 18952 7162 18964
rect 9950 18952 9956 18964
rect 7156 18924 9956 18952
rect 7156 18912 7162 18924
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10502 18912 10508 18964
rect 10560 18912 10566 18964
rect 18322 18912 18328 18964
rect 18380 18952 18386 18964
rect 18966 18952 18972 18964
rect 18380 18924 18972 18952
rect 18380 18912 18386 18924
rect 18966 18912 18972 18924
rect 19024 18912 19030 18964
rect 19426 18912 19432 18964
rect 19484 18912 19490 18964
rect 19797 18955 19855 18961
rect 19797 18921 19809 18955
rect 19843 18952 19855 18955
rect 20346 18952 20352 18964
rect 19843 18924 20352 18952
rect 19843 18921 19855 18924
rect 19797 18915 19855 18921
rect 20346 18912 20352 18924
rect 20404 18912 20410 18964
rect 21726 18912 21732 18964
rect 21784 18912 21790 18964
rect 21910 18912 21916 18964
rect 21968 18952 21974 18964
rect 23842 18952 23848 18964
rect 21968 18924 23848 18952
rect 21968 18912 21974 18924
rect 23842 18912 23848 18924
rect 23900 18912 23906 18964
rect 9030 18844 9036 18896
rect 9088 18884 9094 18896
rect 9306 18884 9312 18896
rect 9088 18856 9312 18884
rect 9088 18844 9094 18856
rect 9306 18844 9312 18856
rect 9364 18884 9370 18896
rect 23661 18887 23719 18893
rect 9364 18856 11284 18884
rect 9364 18844 9370 18856
rect 7469 18819 7527 18825
rect 7469 18785 7481 18819
rect 7515 18816 7527 18819
rect 10781 18819 10839 18825
rect 10781 18816 10793 18819
rect 7515 18788 10793 18816
rect 7515 18785 7527 18788
rect 7469 18779 7527 18785
rect 10781 18785 10793 18788
rect 10827 18785 10839 18819
rect 10781 18779 10839 18785
rect 10870 18776 10876 18828
rect 10928 18776 10934 18828
rect 11256 18825 11284 18856
rect 23661 18853 23673 18887
rect 23707 18884 23719 18887
rect 24670 18884 24676 18896
rect 23707 18856 24676 18884
rect 23707 18853 23719 18856
rect 23661 18847 23719 18853
rect 24670 18844 24676 18856
rect 24728 18844 24734 18896
rect 11241 18819 11299 18825
rect 11241 18785 11253 18819
rect 11287 18785 11299 18819
rect 11241 18779 11299 18785
rect 15105 18819 15163 18825
rect 15105 18785 15117 18819
rect 15151 18816 15163 18819
rect 15838 18816 15844 18828
rect 15151 18788 15844 18816
rect 15151 18785 15163 18788
rect 15105 18779 15163 18785
rect 15838 18776 15844 18788
rect 15896 18776 15902 18828
rect 19337 18819 19395 18825
rect 19337 18785 19349 18819
rect 19383 18816 19395 18819
rect 20254 18816 20260 18828
rect 19383 18788 20260 18816
rect 19383 18785 19395 18788
rect 19337 18779 19395 18785
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 23385 18819 23443 18825
rect 23385 18785 23397 18819
rect 23431 18816 23443 18819
rect 24026 18816 24032 18828
rect 23431 18788 24032 18816
rect 23431 18785 23443 18788
rect 23385 18779 23443 18785
rect 24026 18776 24032 18788
rect 24084 18776 24090 18828
rect 24486 18776 24492 18828
rect 24544 18776 24550 18828
rect 3786 18708 3792 18760
rect 3844 18748 3850 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3844 18720 4077 18748
rect 3844 18708 3850 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18748 4307 18751
rect 4614 18748 4620 18760
rect 4295 18720 4620 18748
rect 4295 18717 4307 18720
rect 4249 18711 4307 18717
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 5258 18708 5264 18760
rect 5316 18708 5322 18760
rect 7193 18751 7251 18757
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 7558 18748 7564 18760
rect 7239 18720 7564 18748
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 9030 18708 9036 18760
rect 9088 18708 9094 18760
rect 9214 18708 9220 18760
rect 9272 18708 9278 18760
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18717 9459 18751
rect 9401 18711 9459 18717
rect 5534 18689 5540 18692
rect 5528 18643 5540 18689
rect 5534 18640 5540 18643
rect 5592 18640 5598 18692
rect 6914 18640 6920 18692
rect 6972 18640 6978 18692
rect 7285 18683 7343 18689
rect 7285 18680 7297 18683
rect 7024 18652 7297 18680
rect 4433 18615 4491 18621
rect 4433 18581 4445 18615
rect 4479 18612 4491 18615
rect 4798 18612 4804 18624
rect 4479 18584 4804 18612
rect 4479 18581 4491 18584
rect 4433 18575 4491 18581
rect 4798 18572 4804 18584
rect 4856 18572 4862 18624
rect 6638 18572 6644 18624
rect 6696 18572 6702 18624
rect 6730 18572 6736 18624
rect 6788 18612 6794 18624
rect 7024 18612 7052 18652
rect 7285 18649 7297 18652
rect 7331 18649 7343 18683
rect 7285 18643 7343 18649
rect 7745 18683 7803 18689
rect 7745 18649 7757 18683
rect 7791 18649 7803 18683
rect 7745 18643 7803 18649
rect 6788 18584 7052 18612
rect 6788 18572 6794 18584
rect 7098 18572 7104 18624
rect 7156 18572 7162 18624
rect 7760 18612 7788 18643
rect 7834 18640 7840 18692
rect 7892 18680 7898 18692
rect 9309 18683 9367 18689
rect 9309 18680 9321 18683
rect 7892 18652 9321 18680
rect 7892 18640 7898 18652
rect 9309 18649 9321 18652
rect 9355 18649 9367 18683
rect 9416 18680 9444 18711
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9640 18720 9873 18748
rect 9640 18708 9646 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 10008 18720 11161 18748
rect 10008 18708 10014 18720
rect 11149 18717 11161 18720
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 15979 18720 17601 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 17589 18717 17601 18720
rect 17635 18748 17647 18751
rect 18138 18748 18144 18760
rect 17635 18720 18144 18748
rect 17635 18717 17647 18720
rect 17589 18711 17647 18717
rect 18138 18708 18144 18720
rect 18196 18748 18202 18760
rect 18598 18748 18604 18760
rect 18196 18720 18604 18748
rect 18196 18708 18202 18720
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 11425 18683 11483 18689
rect 11425 18680 11437 18683
rect 9416 18652 11437 18680
rect 9309 18643 9367 18649
rect 11425 18649 11437 18652
rect 11471 18649 11483 18683
rect 11425 18643 11483 18649
rect 15657 18683 15715 18689
rect 15657 18649 15669 18683
rect 15703 18680 15715 18683
rect 16178 18683 16236 18689
rect 16178 18680 16190 18683
rect 15703 18652 16190 18680
rect 15703 18649 15715 18652
rect 15657 18643 15715 18649
rect 16178 18649 16190 18652
rect 16224 18649 16236 18683
rect 16178 18643 16236 18649
rect 17402 18640 17408 18692
rect 17460 18680 17466 18692
rect 17834 18683 17892 18689
rect 17834 18680 17846 18683
rect 17460 18652 17846 18680
rect 17460 18640 17466 18652
rect 17834 18649 17846 18652
rect 17880 18649 17892 18683
rect 17834 18643 17892 18649
rect 9398 18612 9404 18624
rect 7760 18584 9404 18612
rect 9398 18572 9404 18584
rect 9456 18572 9462 18624
rect 9585 18615 9643 18621
rect 9585 18581 9597 18615
rect 9631 18612 9643 18615
rect 10686 18612 10692 18624
rect 9631 18584 10692 18612
rect 9631 18581 9643 18584
rect 9585 18575 9643 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 10962 18572 10968 18624
rect 11020 18572 11026 18624
rect 17310 18572 17316 18624
rect 17368 18572 17374 18624
rect 19628 18612 19656 18711
rect 20162 18708 20168 18760
rect 20220 18748 20226 18760
rect 20349 18751 20407 18757
rect 20349 18748 20361 18751
rect 20220 18720 20361 18748
rect 20220 18708 20226 18720
rect 20349 18717 20361 18720
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 23106 18708 23112 18760
rect 23164 18757 23170 18760
rect 23164 18748 23176 18757
rect 23164 18720 23209 18748
rect 23164 18711 23176 18720
rect 23164 18708 23170 18711
rect 23658 18708 23664 18760
rect 23716 18708 23722 18760
rect 23937 18751 23995 18757
rect 23937 18717 23949 18751
rect 23983 18717 23995 18751
rect 23937 18711 23995 18717
rect 20616 18683 20674 18689
rect 20616 18649 20628 18683
rect 20662 18680 20674 18683
rect 20806 18680 20812 18692
rect 20662 18652 20812 18680
rect 20662 18649 20674 18652
rect 20616 18643 20674 18649
rect 20806 18640 20812 18652
rect 20864 18640 20870 18692
rect 23952 18680 23980 18711
rect 24854 18680 24860 18692
rect 23952 18652 24860 18680
rect 24854 18640 24860 18652
rect 24912 18680 24918 18692
rect 25133 18683 25191 18689
rect 25133 18680 25145 18683
rect 24912 18652 25145 18680
rect 24912 18640 24918 18652
rect 25133 18649 25145 18652
rect 25179 18649 25191 18683
rect 25133 18643 25191 18649
rect 20714 18612 20720 18624
rect 19628 18584 20720 18612
rect 20714 18572 20720 18584
rect 20772 18572 20778 18624
rect 21910 18572 21916 18624
rect 21968 18612 21974 18624
rect 22005 18615 22063 18621
rect 22005 18612 22017 18615
rect 21968 18584 22017 18612
rect 21968 18572 21974 18584
rect 22005 18581 22017 18584
rect 22051 18581 22063 18615
rect 22005 18575 22063 18581
rect 23842 18572 23848 18624
rect 23900 18572 23906 18624
rect 1104 18522 28888 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 28888 18522
rect 1104 18448 28888 18470
rect 3786 18368 3792 18420
rect 3844 18368 3850 18420
rect 6089 18411 6147 18417
rect 6089 18377 6101 18411
rect 6135 18408 6147 18411
rect 7098 18408 7104 18420
rect 6135 18380 7104 18408
rect 6135 18377 6147 18380
rect 6089 18371 6147 18377
rect 7098 18368 7104 18380
rect 7156 18368 7162 18420
rect 7834 18368 7840 18420
rect 7892 18368 7898 18420
rect 9398 18368 9404 18420
rect 9456 18368 9462 18420
rect 15650 18411 15708 18417
rect 15650 18377 15662 18411
rect 15696 18408 15708 18411
rect 15696 18380 17356 18408
rect 15696 18377 15708 18380
rect 15650 18371 15708 18377
rect 5258 18340 5264 18352
rect 4724 18312 5264 18340
rect 4724 18281 4752 18312
rect 5258 18300 5264 18312
rect 5316 18300 5322 18352
rect 9582 18340 9588 18352
rect 6656 18312 9588 18340
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18241 4767 18275
rect 4709 18235 4767 18241
rect 4976 18275 5034 18281
rect 4976 18241 4988 18275
rect 5022 18272 5034 18275
rect 5442 18272 5448 18284
rect 5022 18244 5448 18272
rect 5022 18241 5034 18244
rect 4976 18235 5034 18241
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 6656 18281 6684 18312
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 16206 18349 16212 18352
rect 16193 18343 16212 18349
rect 16193 18309 16205 18343
rect 16193 18303 16212 18309
rect 16206 18300 16212 18303
rect 16264 18300 16270 18352
rect 16390 18300 16396 18352
rect 16448 18300 16454 18352
rect 16666 18300 16672 18352
rect 16724 18340 16730 18352
rect 16761 18343 16819 18349
rect 16761 18340 16773 18343
rect 16724 18312 16773 18340
rect 16724 18300 16730 18312
rect 16761 18309 16773 18312
rect 16807 18309 16819 18343
rect 16761 18303 16819 18309
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18241 6699 18275
rect 6641 18235 6699 18241
rect 6730 18232 6736 18284
rect 6788 18232 6794 18284
rect 6917 18275 6975 18281
rect 6917 18241 6929 18275
rect 6963 18272 6975 18275
rect 7006 18272 7012 18284
rect 6963 18244 7012 18272
rect 6963 18241 6975 18244
rect 6917 18235 6975 18241
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18272 8171 18275
rect 11057 18275 11115 18281
rect 11057 18272 11069 18275
rect 8159 18244 11069 18272
rect 8159 18241 8171 18244
rect 8113 18235 8171 18241
rect 11057 18241 11069 18244
rect 11103 18272 11115 18275
rect 11330 18272 11336 18284
rect 11103 18244 11336 18272
rect 11103 18241 11115 18244
rect 11057 18235 11115 18241
rect 11330 18232 11336 18244
rect 11388 18272 11394 18284
rect 15473 18275 15531 18281
rect 11388 18244 12434 18272
rect 11388 18232 11394 18244
rect 4433 18207 4491 18213
rect 4433 18173 4445 18207
rect 4479 18173 4491 18207
rect 4433 18167 4491 18173
rect 7285 18207 7343 18213
rect 7285 18173 7297 18207
rect 7331 18204 7343 18207
rect 8202 18204 8208 18216
rect 7331 18176 8208 18204
rect 7331 18173 7343 18176
rect 7285 18167 7343 18173
rect 4448 18136 4476 18167
rect 8202 18164 8208 18176
rect 8260 18164 8266 18216
rect 10686 18164 10692 18216
rect 10744 18164 10750 18216
rect 12158 18164 12164 18216
rect 12216 18164 12222 18216
rect 4706 18136 4712 18148
rect 4448 18108 4712 18136
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 6457 18139 6515 18145
rect 6457 18105 6469 18139
rect 6503 18136 6515 18139
rect 10042 18136 10048 18148
rect 6503 18108 10048 18136
rect 6503 18105 6515 18108
rect 6457 18099 6515 18105
rect 10042 18096 10048 18108
rect 10100 18096 10106 18148
rect 12406 18136 12434 18244
rect 15473 18241 15485 18275
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18272 15623 18275
rect 15654 18272 15660 18284
rect 15611 18244 15660 18272
rect 15611 18241 15623 18244
rect 15565 18235 15623 18241
rect 15378 18164 15384 18216
rect 15436 18204 15442 18216
rect 15488 18204 15516 18235
rect 15654 18232 15660 18244
rect 15712 18232 15718 18284
rect 17328 18281 17356 18380
rect 20806 18368 20812 18420
rect 20864 18368 20870 18420
rect 22370 18368 22376 18420
rect 22428 18368 22434 18420
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18272 15807 18275
rect 17313 18275 17371 18281
rect 15795 18244 16804 18272
rect 15795 18241 15807 18244
rect 15749 18235 15807 18241
rect 16776 18216 16804 18244
rect 17313 18241 17325 18275
rect 17359 18241 17371 18275
rect 17313 18235 17371 18241
rect 18598 18232 18604 18284
rect 18656 18272 18662 18284
rect 20162 18272 20168 18284
rect 18656 18244 20168 18272
rect 18656 18232 18662 18244
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20990 18232 20996 18284
rect 21048 18232 21054 18284
rect 21177 18275 21235 18281
rect 21177 18241 21189 18275
rect 21223 18272 21235 18275
rect 21358 18272 21364 18284
rect 21223 18244 21364 18272
rect 21223 18241 21235 18244
rect 21177 18235 21235 18241
rect 21358 18232 21364 18244
rect 21416 18232 21422 18284
rect 21818 18232 21824 18284
rect 21876 18272 21882 18284
rect 21913 18275 21971 18281
rect 21913 18272 21925 18275
rect 21876 18244 21925 18272
rect 21876 18232 21882 18244
rect 21913 18241 21925 18244
rect 21959 18241 21971 18275
rect 21913 18235 21971 18241
rect 22002 18232 22008 18284
rect 22060 18232 22066 18284
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18272 22247 18275
rect 22554 18272 22560 18284
rect 22235 18244 22560 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 23773 18275 23831 18281
rect 23773 18241 23785 18275
rect 23819 18272 23831 18275
rect 23934 18272 23940 18284
rect 23819 18244 23940 18272
rect 23819 18241 23831 18244
rect 23773 18235 23831 18241
rect 23934 18232 23940 18244
rect 23992 18232 23998 18284
rect 24026 18232 24032 18284
rect 24084 18232 24090 18284
rect 16298 18204 16304 18216
rect 15436 18176 16304 18204
rect 15436 18164 15442 18176
rect 16298 18164 16304 18176
rect 16356 18164 16362 18216
rect 16758 18164 16764 18216
rect 16816 18164 16822 18216
rect 21082 18164 21088 18216
rect 21140 18204 21146 18216
rect 21269 18207 21327 18213
rect 21269 18204 21281 18207
rect 21140 18176 21281 18204
rect 21140 18164 21146 18176
rect 21269 18173 21281 18176
rect 21315 18173 21327 18207
rect 21269 18167 21327 18173
rect 16850 18136 16856 18148
rect 12406 18108 16856 18136
rect 16850 18096 16856 18108
rect 16908 18136 16914 18148
rect 18046 18136 18052 18148
rect 16908 18108 18052 18136
rect 16908 18096 16914 18108
rect 18046 18096 18052 18108
rect 18104 18096 18110 18148
rect 842 18028 848 18080
rect 900 18068 906 18080
rect 1489 18071 1547 18077
rect 1489 18068 1501 18071
rect 900 18040 1501 18068
rect 900 18028 906 18040
rect 1489 18037 1501 18040
rect 1535 18037 1547 18071
rect 1489 18031 1547 18037
rect 6917 18071 6975 18077
rect 6917 18037 6929 18071
rect 6963 18068 6975 18071
rect 7558 18068 7564 18080
rect 6963 18040 7564 18068
rect 6963 18037 6975 18040
rect 6917 18031 6975 18037
rect 7558 18028 7564 18040
rect 7616 18028 7622 18080
rect 10134 18028 10140 18080
rect 10192 18028 10198 18080
rect 11609 18071 11667 18077
rect 11609 18037 11621 18071
rect 11655 18068 11667 18071
rect 11790 18068 11796 18080
rect 11655 18040 11796 18068
rect 11655 18037 11667 18040
rect 11609 18031 11667 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 16022 18028 16028 18080
rect 16080 18028 16086 18080
rect 16209 18071 16267 18077
rect 16209 18037 16221 18071
rect 16255 18068 16267 18071
rect 16758 18068 16764 18080
rect 16255 18040 16764 18068
rect 16255 18037 16267 18040
rect 16209 18031 16267 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 22646 18028 22652 18080
rect 22704 18028 22710 18080
rect 1104 17978 28888 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 28888 17978
rect 1104 17904 28888 17926
rect 5997 17867 6055 17873
rect 5997 17833 6009 17867
rect 6043 17864 6055 17867
rect 7190 17864 7196 17876
rect 6043 17836 7196 17864
rect 6043 17833 6055 17836
rect 5997 17827 6055 17833
rect 7190 17824 7196 17836
rect 7248 17824 7254 17876
rect 8202 17824 8208 17876
rect 8260 17824 8266 17876
rect 9490 17824 9496 17876
rect 9548 17864 9554 17876
rect 10594 17864 10600 17876
rect 9548 17836 10600 17864
rect 9548 17824 9554 17836
rect 10594 17824 10600 17836
rect 10652 17864 10658 17876
rect 11606 17864 11612 17876
rect 10652 17836 11612 17864
rect 10652 17824 10658 17836
rect 11606 17824 11612 17836
rect 11664 17864 11670 17876
rect 11701 17867 11759 17873
rect 11701 17864 11713 17867
rect 11664 17836 11713 17864
rect 11664 17824 11670 17836
rect 11701 17833 11713 17836
rect 11747 17833 11759 17867
rect 11701 17827 11759 17833
rect 16758 17824 16764 17876
rect 16816 17824 16822 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 20993 17867 21051 17873
rect 20993 17864 21005 17867
rect 20772 17836 21005 17864
rect 20772 17824 20778 17836
rect 20993 17833 21005 17836
rect 21039 17833 21051 17867
rect 20993 17827 21051 17833
rect 23934 17824 23940 17876
rect 23992 17864 23998 17876
rect 24489 17867 24547 17873
rect 24489 17864 24501 17867
rect 23992 17836 24501 17864
rect 23992 17824 23998 17836
rect 24489 17833 24501 17836
rect 24535 17833 24547 17867
rect 24489 17827 24547 17833
rect 24854 17824 24860 17876
rect 24912 17824 24918 17876
rect 4614 17756 4620 17808
rect 4672 17756 4678 17808
rect 11333 17799 11391 17805
rect 11333 17765 11345 17799
rect 11379 17796 11391 17799
rect 12434 17796 12440 17808
rect 11379 17768 12440 17796
rect 11379 17765 11391 17768
rect 11333 17759 11391 17765
rect 12434 17756 12440 17768
rect 12492 17756 12498 17808
rect 19521 17799 19579 17805
rect 19521 17765 19533 17799
rect 19567 17796 19579 17799
rect 20898 17796 20904 17808
rect 19567 17768 20904 17796
rect 19567 17765 19579 17768
rect 19521 17759 19579 17765
rect 20898 17756 20904 17768
rect 20956 17756 20962 17808
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 4632 17728 4660 17756
rect 3007 17700 4660 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9953 17731 10011 17737
rect 9953 17728 9965 17731
rect 9456 17700 9965 17728
rect 9456 17688 9462 17700
rect 9953 17697 9965 17700
rect 9999 17697 10011 17731
rect 17310 17728 17316 17740
rect 9953 17691 10011 17697
rect 16316 17700 17316 17728
rect 3142 17620 3148 17672
rect 3200 17620 3206 17672
rect 4617 17663 4675 17669
rect 4617 17629 4629 17663
rect 4663 17629 4675 17663
rect 4617 17623 4675 17629
rect 4884 17663 4942 17669
rect 4884 17629 4896 17663
rect 4930 17629 4942 17663
rect 4884 17623 4942 17629
rect 4632 17536 4660 17623
rect 4798 17552 4804 17604
rect 4856 17592 4862 17604
rect 4908 17592 4936 17623
rect 5258 17620 5264 17672
rect 5316 17660 5322 17672
rect 6825 17663 6883 17669
rect 6825 17660 6837 17663
rect 5316 17632 6837 17660
rect 5316 17620 5322 17632
rect 6825 17629 6837 17632
rect 6871 17660 6883 17663
rect 8018 17660 8024 17672
rect 6871 17632 8024 17660
rect 6871 17629 6883 17632
rect 6825 17623 6883 17629
rect 8018 17620 8024 17632
rect 8076 17620 8082 17672
rect 9306 17620 9312 17672
rect 9364 17620 9370 17672
rect 9490 17620 9496 17672
rect 9548 17620 9554 17672
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17660 9735 17663
rect 11790 17660 11796 17672
rect 9723 17632 11796 17660
rect 9723 17629 9735 17632
rect 9677 17623 9735 17629
rect 11790 17620 11796 17632
rect 11848 17620 11854 17672
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 12161 17663 12219 17669
rect 12161 17660 12173 17663
rect 11940 17632 12173 17660
rect 11940 17620 11946 17632
rect 12161 17629 12173 17632
rect 12207 17660 12219 17663
rect 12250 17660 12256 17672
rect 12207 17632 12256 17660
rect 12207 17629 12219 17632
rect 12161 17623 12219 17629
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 14734 17620 14740 17672
rect 14792 17660 14798 17672
rect 15013 17663 15071 17669
rect 15013 17660 15025 17663
rect 14792 17632 15025 17660
rect 14792 17620 14798 17632
rect 15013 17629 15025 17632
rect 15059 17629 15071 17663
rect 15013 17623 15071 17629
rect 15105 17663 15163 17669
rect 15105 17629 15117 17663
rect 15151 17660 15163 17663
rect 15194 17660 15200 17672
rect 15151 17632 15200 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 15286 17620 15292 17672
rect 15344 17620 15350 17672
rect 15378 17620 15384 17672
rect 15436 17620 15442 17672
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 16316 17669 16344 17700
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 19337 17731 19395 17737
rect 19337 17728 19349 17731
rect 17880 17700 19349 17728
rect 15933 17663 15991 17669
rect 15933 17660 15945 17663
rect 15896 17632 15945 17660
rect 15896 17620 15902 17632
rect 15933 17629 15945 17632
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17629 16359 17663
rect 17218 17660 17224 17672
rect 16301 17623 16359 17629
rect 16408 17632 17224 17660
rect 4856 17564 4936 17592
rect 4856 17552 4862 17564
rect 3329 17527 3387 17533
rect 3329 17493 3341 17527
rect 3375 17524 3387 17527
rect 3418 17524 3424 17536
rect 3375 17496 3424 17524
rect 3375 17493 3387 17496
rect 3329 17487 3387 17493
rect 3418 17484 3424 17496
rect 3476 17484 3482 17536
rect 4614 17484 4620 17536
rect 4672 17524 4678 17536
rect 5276 17524 5304 17620
rect 6086 17552 6092 17604
rect 6144 17592 6150 17604
rect 7070 17595 7128 17601
rect 7070 17592 7082 17595
rect 6144 17564 7082 17592
rect 6144 17552 6150 17564
rect 7070 17561 7082 17564
rect 7116 17561 7128 17595
rect 9324 17592 9352 17620
rect 10198 17595 10256 17601
rect 10198 17592 10210 17595
rect 9324 17564 10210 17592
rect 7070 17555 7128 17561
rect 10198 17561 10210 17564
rect 10244 17561 10256 17595
rect 10198 17555 10256 17561
rect 15565 17595 15623 17601
rect 15565 17561 15577 17595
rect 15611 17592 15623 17595
rect 16117 17595 16175 17601
rect 16117 17592 16129 17595
rect 15611 17564 16129 17592
rect 15611 17561 15623 17564
rect 15565 17555 15623 17561
rect 16117 17561 16129 17564
rect 16163 17561 16175 17595
rect 16117 17555 16175 17561
rect 16209 17595 16267 17601
rect 16209 17561 16221 17595
rect 16255 17592 16267 17595
rect 16408 17592 16436 17632
rect 17218 17620 17224 17632
rect 17276 17620 17282 17672
rect 17880 17669 17908 17700
rect 19337 17697 19349 17700
rect 19383 17697 19395 17731
rect 19337 17691 19395 17697
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 20622 17728 20628 17740
rect 19843 17700 20628 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 20622 17688 20628 17700
rect 20680 17688 20686 17740
rect 20916 17700 21772 17728
rect 17865 17663 17923 17669
rect 17865 17629 17877 17663
rect 17911 17629 17923 17663
rect 17865 17623 17923 17629
rect 17954 17620 17960 17672
rect 18012 17620 18018 17672
rect 18322 17620 18328 17672
rect 18380 17669 18386 17672
rect 18380 17660 18388 17669
rect 20165 17663 20223 17669
rect 20165 17660 20177 17663
rect 18380 17632 18425 17660
rect 18524 17632 20177 17660
rect 18380 17623 18388 17632
rect 18380 17620 18386 17623
rect 18141 17595 18199 17601
rect 18141 17592 18153 17595
rect 16255 17564 16436 17592
rect 16500 17564 18153 17592
rect 16255 17561 16267 17564
rect 16209 17555 16267 17561
rect 4672 17496 5304 17524
rect 4672 17484 4678 17496
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 9490 17524 9496 17536
rect 5960 17496 9496 17524
rect 5960 17484 5966 17496
rect 9490 17484 9496 17496
rect 9548 17484 9554 17536
rect 16500 17533 16528 17564
rect 18141 17561 18153 17564
rect 18187 17561 18199 17595
rect 18141 17555 18199 17561
rect 18230 17552 18236 17604
rect 18288 17552 18294 17604
rect 18524 17533 18552 17632
rect 20165 17629 20177 17632
rect 20211 17629 20223 17663
rect 20165 17623 20223 17629
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17660 20591 17663
rect 20916 17660 20944 17700
rect 21744 17672 21772 17700
rect 22646 17688 22652 17740
rect 22704 17728 22710 17740
rect 23293 17731 23351 17737
rect 23293 17728 23305 17731
rect 22704 17700 23305 17728
rect 22704 17688 22710 17700
rect 23293 17697 23305 17700
rect 23339 17697 23351 17731
rect 23293 17691 23351 17697
rect 23658 17688 23664 17740
rect 23716 17728 23722 17740
rect 23934 17728 23940 17740
rect 23716 17700 23940 17728
rect 23716 17688 23722 17700
rect 23934 17688 23940 17700
rect 23992 17688 23998 17740
rect 20579 17632 20944 17660
rect 20993 17663 21051 17669
rect 20579 17629 20591 17632
rect 20533 17623 20591 17629
rect 20993 17629 21005 17663
rect 21039 17660 21051 17663
rect 21082 17660 21088 17672
rect 21039 17632 21088 17660
rect 21039 17629 21051 17632
rect 20993 17623 21051 17629
rect 21082 17620 21088 17632
rect 21140 17620 21146 17672
rect 21177 17663 21235 17669
rect 21177 17629 21189 17663
rect 21223 17660 21235 17663
rect 21450 17660 21456 17672
rect 21223 17632 21456 17660
rect 21223 17629 21235 17632
rect 21177 17623 21235 17629
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 21545 17663 21603 17669
rect 21545 17629 21557 17663
rect 21591 17629 21603 17663
rect 21545 17623 21603 17629
rect 20346 17552 20352 17604
rect 20404 17552 20410 17604
rect 20441 17595 20499 17601
rect 20441 17561 20453 17595
rect 20487 17561 20499 17595
rect 21560 17592 21588 17623
rect 21726 17620 21732 17672
rect 21784 17620 21790 17672
rect 21818 17620 21824 17672
rect 21876 17620 21882 17672
rect 21910 17620 21916 17672
rect 21968 17620 21974 17672
rect 22097 17663 22155 17669
rect 22097 17629 22109 17663
rect 22143 17660 22155 17663
rect 22186 17660 22192 17672
rect 22143 17632 22192 17660
rect 22143 17629 22155 17632
rect 22097 17623 22155 17629
rect 22186 17620 22192 17632
rect 22244 17620 22250 17672
rect 24670 17620 24676 17672
rect 24728 17620 24734 17672
rect 24949 17663 25007 17669
rect 24949 17629 24961 17663
rect 24995 17629 25007 17663
rect 24949 17623 25007 17629
rect 24964 17592 24992 17623
rect 20441 17555 20499 17561
rect 20916 17564 21588 17592
rect 23952 17564 24992 17592
rect 16485 17527 16543 17533
rect 16485 17493 16497 17527
rect 16531 17493 16543 17527
rect 16485 17487 16543 17493
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17493 18567 17527
rect 20456 17524 20484 17555
rect 20530 17524 20536 17536
rect 20456 17496 20536 17524
rect 18509 17487 18567 17493
rect 20530 17484 20536 17496
rect 20588 17484 20594 17536
rect 20717 17527 20775 17533
rect 20717 17493 20729 17527
rect 20763 17524 20775 17527
rect 20916 17524 20944 17564
rect 20763 17496 20944 17524
rect 22281 17527 22339 17533
rect 20763 17493 20775 17496
rect 20717 17487 20775 17493
rect 22281 17493 22293 17527
rect 22327 17524 22339 17527
rect 23106 17524 23112 17536
rect 22327 17496 23112 17524
rect 22327 17493 22339 17496
rect 22281 17487 22339 17493
rect 23106 17484 23112 17496
rect 23164 17484 23170 17536
rect 23474 17484 23480 17536
rect 23532 17524 23538 17536
rect 23842 17524 23848 17536
rect 23532 17496 23848 17524
rect 23532 17484 23538 17496
rect 23842 17484 23848 17496
rect 23900 17524 23906 17536
rect 23952 17533 23980 17564
rect 23937 17527 23995 17533
rect 23937 17524 23949 17527
rect 23900 17496 23949 17524
rect 23900 17484 23906 17496
rect 23937 17493 23949 17496
rect 23983 17493 23995 17527
rect 23937 17487 23995 17493
rect 1104 17434 28888 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 28888 17434
rect 1104 17360 28888 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 3142 17320 3148 17332
rect 1719 17292 3148 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 3142 17280 3148 17292
rect 3200 17280 3206 17332
rect 5445 17323 5503 17329
rect 5445 17289 5457 17323
rect 5491 17320 5503 17323
rect 5534 17320 5540 17332
rect 5491 17292 5540 17320
rect 5491 17289 5503 17292
rect 5445 17283 5503 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 6086 17280 6092 17332
rect 6144 17280 6150 17332
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 7282 17320 7288 17332
rect 6972 17292 7288 17320
rect 6972 17280 6978 17292
rect 7282 17280 7288 17292
rect 7340 17320 7346 17332
rect 7377 17323 7435 17329
rect 7377 17320 7389 17323
rect 7340 17292 7389 17320
rect 7340 17280 7346 17292
rect 7377 17289 7389 17292
rect 7423 17289 7435 17323
rect 7377 17283 7435 17289
rect 9493 17323 9551 17329
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 9582 17320 9588 17332
rect 9539 17292 9588 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 11149 17323 11207 17329
rect 11149 17289 11161 17323
rect 11195 17320 11207 17323
rect 11698 17320 11704 17332
rect 11195 17292 11704 17320
rect 11195 17289 11207 17292
rect 11149 17283 11207 17289
rect 11698 17280 11704 17292
rect 11756 17320 11762 17332
rect 12158 17320 12164 17332
rect 11756 17292 12164 17320
rect 11756 17280 11762 17292
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 15838 17280 15844 17332
rect 15896 17280 15902 17332
rect 17589 17323 17647 17329
rect 17589 17289 17601 17323
rect 17635 17320 17647 17323
rect 17954 17320 17960 17332
rect 17635 17292 17960 17320
rect 17635 17289 17647 17292
rect 17589 17283 17647 17289
rect 17954 17280 17960 17292
rect 18012 17280 18018 17332
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 18104 17292 18460 17320
rect 18104 17280 18110 17292
rect 4614 17252 4620 17264
rect 3344 17224 4620 17252
rect 1302 17144 1308 17196
rect 1360 17184 1366 17196
rect 3344 17193 3372 17224
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 6932 17252 6960 17280
rect 5828 17224 6960 17252
rect 1489 17187 1547 17193
rect 1489 17184 1501 17187
rect 1360 17156 1501 17184
rect 1360 17144 1366 17156
rect 1489 17153 1501 17156
rect 1535 17184 1547 17187
rect 1949 17187 2007 17193
rect 1949 17184 1961 17187
rect 1535 17156 1961 17184
rect 1535 17153 1547 17156
rect 1489 17147 1547 17153
rect 1949 17153 1961 17156
rect 1995 17153 2007 17187
rect 1949 17147 2007 17153
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17153 3387 17187
rect 3329 17147 3387 17153
rect 3418 17144 3424 17196
rect 3476 17184 3482 17196
rect 5828 17193 5856 17224
rect 8018 17212 8024 17264
rect 8076 17252 8082 17264
rect 10036 17255 10094 17261
rect 8076 17224 9444 17252
rect 8076 17212 8082 17224
rect 3585 17187 3643 17193
rect 3585 17184 3597 17187
rect 3476 17156 3597 17184
rect 3476 17144 3482 17156
rect 3585 17153 3597 17156
rect 3631 17153 3643 17187
rect 3585 17147 3643 17153
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17184 5319 17187
rect 5813 17187 5871 17193
rect 5307 17156 5764 17184
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17116 5135 17119
rect 5626 17116 5632 17128
rect 5123 17088 5632 17116
rect 5123 17085 5135 17088
rect 5077 17079 5135 17085
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 5736 17116 5764 17156
rect 5813 17153 5825 17187
rect 5859 17153 5871 17187
rect 5813 17147 5871 17153
rect 5902 17144 5908 17196
rect 5960 17144 5966 17196
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 6696 17156 6745 17184
rect 6696 17144 6702 17156
rect 6733 17153 6745 17156
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 5920 17116 5948 17144
rect 5736 17088 5948 17116
rect 8036 17116 8064 17212
rect 9416 17196 9444 17224
rect 10036 17221 10048 17255
rect 10082 17252 10094 17255
rect 10134 17252 10140 17264
rect 10082 17224 10140 17252
rect 10082 17221 10094 17224
rect 10036 17215 10094 17221
rect 10134 17212 10140 17224
rect 10192 17212 10198 17264
rect 15378 17212 15384 17264
rect 15436 17252 15442 17264
rect 15473 17255 15531 17261
rect 15473 17252 15485 17255
rect 15436 17224 15485 17252
rect 15436 17212 15442 17224
rect 15473 17221 15485 17224
rect 15519 17221 15531 17255
rect 18230 17252 18236 17264
rect 15473 17215 15531 17221
rect 17052 17224 18236 17252
rect 8202 17144 8208 17196
rect 8260 17184 8266 17196
rect 8369 17187 8427 17193
rect 8369 17184 8381 17187
rect 8260 17156 8381 17184
rect 8260 17144 8266 17156
rect 8369 17153 8381 17156
rect 8415 17153 8427 17187
rect 8369 17147 8427 17153
rect 9398 17144 9404 17196
rect 9456 17184 9462 17196
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 9456 17156 9781 17184
rect 9456 17144 9462 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 12250 17144 12256 17196
rect 12308 17144 12314 17196
rect 12434 17144 12440 17196
rect 12492 17144 12498 17196
rect 15286 17144 15292 17196
rect 15344 17184 15350 17196
rect 17052 17193 17080 17224
rect 18230 17212 18236 17224
rect 18288 17212 18294 17264
rect 18432 17261 18460 17292
rect 20346 17280 20352 17332
rect 20404 17320 20410 17332
rect 20441 17323 20499 17329
rect 20441 17320 20453 17323
rect 20404 17292 20453 17320
rect 20404 17280 20410 17292
rect 20441 17289 20453 17292
rect 20487 17289 20499 17323
rect 20441 17283 20499 17289
rect 20530 17280 20536 17332
rect 20588 17320 20594 17332
rect 21266 17320 21272 17332
rect 20588 17292 21272 17320
rect 20588 17280 20594 17292
rect 21266 17280 21272 17292
rect 21324 17320 21330 17332
rect 21818 17320 21824 17332
rect 21324 17292 21824 17320
rect 21324 17280 21330 17292
rect 21818 17280 21824 17292
rect 21876 17280 21882 17332
rect 18417 17255 18475 17261
rect 18417 17221 18429 17255
rect 18463 17221 18475 17255
rect 18417 17215 18475 17221
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 15344 17156 15669 17184
rect 15344 17144 15350 17156
rect 15657 17153 15669 17156
rect 15703 17153 15715 17187
rect 15657 17147 15715 17153
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17218 17144 17224 17196
rect 17276 17184 17282 17196
rect 17313 17187 17371 17193
rect 17313 17184 17325 17187
rect 17276 17156 17325 17184
rect 17276 17144 17282 17156
rect 17313 17153 17325 17156
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 17402 17144 17408 17196
rect 17460 17144 17466 17196
rect 20622 17144 20628 17196
rect 20680 17193 20686 17196
rect 20680 17187 20713 17193
rect 20701 17153 20713 17187
rect 20680 17147 20713 17153
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17184 20867 17187
rect 20898 17184 20904 17196
rect 20855 17156 20904 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 20680 17144 20686 17147
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 21910 17144 21916 17196
rect 21968 17184 21974 17196
rect 22373 17187 22431 17193
rect 22373 17184 22385 17187
rect 21968 17156 22385 17184
rect 21968 17144 21974 17156
rect 22373 17153 22385 17156
rect 22419 17153 22431 17187
rect 22373 17147 22431 17153
rect 22557 17187 22615 17193
rect 22557 17153 22569 17187
rect 22603 17184 22615 17187
rect 23017 17187 23075 17193
rect 23017 17184 23029 17187
rect 22603 17156 23029 17184
rect 22603 17153 22615 17156
rect 22557 17147 22615 17153
rect 23017 17153 23029 17156
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 23106 17144 23112 17196
rect 23164 17144 23170 17196
rect 23385 17187 23443 17193
rect 23385 17153 23397 17187
rect 23431 17184 23443 17187
rect 23658 17184 23664 17196
rect 23431 17156 23664 17184
rect 23431 17153 23443 17156
rect 23385 17147 23443 17153
rect 23658 17144 23664 17156
rect 23716 17144 23722 17196
rect 27249 17187 27307 17193
rect 27249 17153 27261 17187
rect 27295 17184 27307 17187
rect 27522 17184 27528 17196
rect 27295 17156 27528 17184
rect 27295 17153 27307 17156
rect 27249 17147 27307 17153
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 8036 17088 8125 17116
rect 8113 17085 8125 17088
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17116 17187 17119
rect 18322 17116 18328 17128
rect 17175 17088 18328 17116
rect 17175 17085 17187 17088
rect 17129 17079 17187 17085
rect 18322 17076 18328 17088
rect 18380 17076 18386 17128
rect 20162 17076 20168 17128
rect 20220 17076 20226 17128
rect 22186 17076 22192 17128
rect 22244 17076 22250 17128
rect 24302 17076 24308 17128
rect 24360 17076 24366 17128
rect 28258 17076 28264 17128
rect 28316 17076 28322 17128
rect 4706 16940 4712 16992
rect 4764 16940 4770 16992
rect 12345 16983 12403 16989
rect 12345 16949 12357 16983
rect 12391 16980 12403 16983
rect 13262 16980 13268 16992
rect 12391 16952 13268 16980
rect 12391 16949 12403 16952
rect 12345 16943 12403 16949
rect 13262 16940 13268 16952
rect 13320 16940 13326 16992
rect 22830 16940 22836 16992
rect 22888 16940 22894 16992
rect 23293 16983 23351 16989
rect 23293 16949 23305 16983
rect 23339 16980 23351 16983
rect 23474 16980 23480 16992
rect 23339 16952 23480 16980
rect 23339 16949 23351 16952
rect 23293 16943 23351 16949
rect 23474 16940 23480 16952
rect 23532 16940 23538 16992
rect 24946 16940 24952 16992
rect 25004 16940 25010 16992
rect 1104 16890 28888 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 28888 16890
rect 1104 16816 28888 16838
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 7469 16779 7527 16785
rect 7469 16776 7481 16779
rect 4764 16748 7481 16776
rect 4764 16736 4770 16748
rect 7469 16745 7481 16748
rect 7515 16745 7527 16779
rect 7469 16739 7527 16745
rect 8113 16779 8171 16785
rect 8113 16745 8125 16779
rect 8159 16776 8171 16779
rect 8202 16776 8208 16788
rect 8159 16748 8208 16776
rect 8159 16745 8171 16748
rect 8113 16739 8171 16745
rect 7484 16708 7512 16739
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 23937 16779 23995 16785
rect 23937 16745 23949 16779
rect 23983 16776 23995 16779
rect 24302 16776 24308 16788
rect 23983 16748 24308 16776
rect 23983 16745 23995 16748
rect 23937 16739 23995 16745
rect 24302 16736 24308 16748
rect 24360 16736 24366 16788
rect 24412 16748 26234 16776
rect 10962 16708 10968 16720
rect 7484 16680 10968 16708
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 11882 16708 11888 16720
rect 11072 16680 11888 16708
rect 6733 16643 6791 16649
rect 6733 16609 6745 16643
rect 6779 16640 6791 16643
rect 7098 16640 7104 16652
rect 6779 16612 7104 16640
rect 6779 16609 6791 16612
rect 6733 16603 6791 16609
rect 7098 16600 7104 16612
rect 7156 16640 7162 16652
rect 7745 16643 7803 16649
rect 7156 16612 7512 16640
rect 7156 16600 7162 16612
rect 5626 16532 5632 16584
rect 5684 16572 5690 16584
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 5684 16544 6101 16572
rect 5684 16532 5690 16544
rect 6089 16541 6101 16544
rect 6135 16541 6147 16575
rect 6089 16535 6147 16541
rect 7190 16532 7196 16584
rect 7248 16532 7254 16584
rect 7282 16532 7288 16584
rect 7340 16532 7346 16584
rect 7484 16581 7512 16612
rect 7745 16609 7757 16643
rect 7791 16640 7803 16643
rect 7834 16640 7840 16652
rect 7791 16612 7840 16640
rect 7791 16609 7803 16612
rect 7745 16603 7803 16609
rect 7834 16600 7840 16612
rect 7892 16600 7898 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 7944 16612 8401 16640
rect 7944 16581 7972 16612
rect 8389 16609 8401 16612
rect 8435 16640 8447 16643
rect 11072 16640 11100 16680
rect 11882 16668 11888 16680
rect 11940 16668 11946 16720
rect 24412 16708 24440 16748
rect 23952 16680 24440 16708
rect 8435 16612 11100 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 11793 16643 11851 16649
rect 11793 16640 11805 16643
rect 11756 16612 11805 16640
rect 11756 16600 11762 16612
rect 11793 16609 11805 16612
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 12526 16600 12532 16652
rect 12584 16600 12590 16652
rect 12636 16612 13308 16640
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16541 7527 16575
rect 7469 16535 7527 16541
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 11882 16532 11888 16584
rect 11940 16572 11946 16584
rect 12161 16575 12219 16581
rect 12161 16572 12173 16575
rect 11940 16544 12173 16572
rect 11940 16532 11946 16544
rect 12161 16541 12173 16544
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12636 16572 12664 16612
rect 13280 16581 13308 16612
rect 22830 16600 22836 16652
rect 22888 16640 22894 16652
rect 23845 16643 23903 16649
rect 23845 16640 23857 16643
rect 22888 16612 23857 16640
rect 22888 16600 22894 16612
rect 23845 16609 23857 16612
rect 23891 16609 23903 16643
rect 23845 16603 23903 16609
rect 23952 16584 23980 16680
rect 24026 16600 24032 16652
rect 24084 16640 24090 16652
rect 24673 16643 24731 16649
rect 24673 16640 24685 16643
rect 24084 16612 24685 16640
rect 24084 16600 24090 16612
rect 24673 16609 24685 16612
rect 24719 16609 24731 16643
rect 26206 16640 26234 16748
rect 27522 16736 27528 16788
rect 27580 16736 27586 16788
rect 26206 16612 27752 16640
rect 24673 16603 24731 16609
rect 12492 16544 12664 16572
rect 12713 16575 12771 16581
rect 12492 16532 12498 16544
rect 12713 16541 12725 16575
rect 12759 16541 12771 16575
rect 12713 16535 12771 16541
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16541 13323 16575
rect 13265 16535 13323 16541
rect 12250 16464 12256 16516
rect 12308 16504 12314 16516
rect 12728 16504 12756 16535
rect 23474 16532 23480 16584
rect 23532 16532 23538 16584
rect 23753 16575 23811 16581
rect 23753 16541 23765 16575
rect 23799 16572 23811 16575
rect 23934 16572 23940 16584
rect 23799 16544 23940 16572
rect 23799 16541 23811 16544
rect 23753 16535 23811 16541
rect 23934 16532 23940 16544
rect 23992 16532 23998 16584
rect 24946 16581 24952 16584
rect 24940 16535 24952 16581
rect 24946 16532 24952 16535
rect 25004 16532 25010 16584
rect 27724 16581 27752 16612
rect 27709 16575 27767 16581
rect 27709 16541 27721 16575
rect 27755 16574 27767 16575
rect 27985 16575 28043 16581
rect 27755 16572 27789 16574
rect 27985 16572 27997 16575
rect 27755 16544 27997 16572
rect 27755 16541 27767 16544
rect 27709 16535 27767 16541
rect 27985 16541 27997 16544
rect 28031 16541 28043 16575
rect 27985 16535 28043 16541
rect 13081 16507 13139 16513
rect 13081 16504 13093 16507
rect 12308 16476 13093 16504
rect 12308 16464 12314 16476
rect 13081 16473 13093 16476
rect 13127 16473 13139 16507
rect 13081 16467 13139 16473
rect 7006 16396 7012 16448
rect 7064 16396 7070 16448
rect 13170 16396 13176 16448
rect 13228 16436 13234 16448
rect 13449 16439 13507 16445
rect 13449 16436 13461 16439
rect 13228 16408 13461 16436
rect 13228 16396 13234 16408
rect 13449 16405 13461 16408
rect 13495 16405 13507 16439
rect 13449 16399 13507 16405
rect 23569 16439 23627 16445
rect 23569 16405 23581 16439
rect 23615 16436 23627 16439
rect 23658 16436 23664 16448
rect 23615 16408 23664 16436
rect 23615 16405 23627 16408
rect 23569 16399 23627 16405
rect 23658 16396 23664 16408
rect 23716 16396 23722 16448
rect 26053 16439 26111 16445
rect 26053 16405 26065 16439
rect 26099 16436 26111 16439
rect 27062 16436 27068 16448
rect 26099 16408 27068 16436
rect 26099 16405 26111 16408
rect 26053 16399 26111 16405
rect 27062 16396 27068 16408
rect 27120 16396 27126 16448
rect 1104 16346 28888 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 28888 16346
rect 1104 16272 28888 16294
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 13630 16232 13636 16244
rect 12584 16204 13636 16232
rect 12584 16192 12590 16204
rect 13630 16192 13636 16204
rect 13688 16232 13694 16244
rect 14001 16235 14059 16241
rect 14001 16232 14013 16235
rect 13688 16204 14013 16232
rect 13688 16192 13694 16204
rect 14001 16201 14013 16204
rect 14047 16201 14059 16235
rect 14001 16195 14059 16201
rect 15286 16164 15292 16176
rect 14200 16136 15292 16164
rect 11790 16056 11796 16108
rect 11848 16056 11854 16108
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 11882 15988 11888 16040
rect 11940 15988 11946 16040
rect 12161 15963 12219 15969
rect 12161 15929 12173 15963
rect 12207 15960 12219 15963
rect 12452 15960 12480 16059
rect 13170 16056 13176 16108
rect 13228 16056 13234 16108
rect 13262 16056 13268 16108
rect 13320 16056 13326 16108
rect 13906 16056 13912 16108
rect 13964 16056 13970 16108
rect 14200 16105 14228 16136
rect 15286 16124 15292 16136
rect 15344 16124 15350 16176
rect 14185 16099 14243 16105
rect 14185 16065 14197 16099
rect 14231 16065 14243 16099
rect 14185 16059 14243 16065
rect 14274 16056 14280 16108
rect 14332 16096 14338 16108
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 14332 16068 14657 16096
rect 14332 16056 14338 16068
rect 14645 16065 14657 16068
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 27062 16056 27068 16108
rect 27120 16056 27126 16108
rect 28258 15988 28264 16040
rect 28316 15988 28322 16040
rect 12207 15932 12480 15960
rect 12713 15963 12771 15969
rect 12207 15929 12219 15932
rect 12161 15923 12219 15929
rect 12713 15929 12725 15963
rect 12759 15929 12771 15963
rect 12713 15923 12771 15929
rect 14369 15963 14427 15969
rect 14369 15929 14381 15963
rect 14415 15960 14427 15963
rect 15746 15960 15752 15972
rect 14415 15932 15752 15960
rect 14415 15929 14427 15932
rect 14369 15923 14427 15929
rect 12728 15892 12756 15923
rect 15746 15920 15752 15932
rect 15804 15920 15810 15972
rect 14458 15892 14464 15904
rect 12728 15864 14464 15892
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 14734 15852 14740 15904
rect 14792 15852 14798 15904
rect 23934 15852 23940 15904
rect 23992 15892 23998 15904
rect 24029 15895 24087 15901
rect 24029 15892 24041 15895
rect 23992 15864 24041 15892
rect 23992 15852 23998 15864
rect 24029 15861 24041 15864
rect 24075 15861 24087 15895
rect 24029 15855 24087 15861
rect 1104 15802 28888 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 28888 15802
rect 1104 15728 28888 15750
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12713 15691 12771 15697
rect 12713 15688 12725 15691
rect 12492 15660 12725 15688
rect 12492 15648 12498 15660
rect 12713 15657 12725 15660
rect 12759 15657 12771 15691
rect 12713 15651 12771 15657
rect 13630 15648 13636 15700
rect 13688 15648 13694 15700
rect 14826 15648 14832 15700
rect 14884 15648 14890 15700
rect 12069 15623 12127 15629
rect 12069 15589 12081 15623
rect 12115 15589 12127 15623
rect 12069 15583 12127 15589
rect 13817 15623 13875 15629
rect 13817 15589 13829 15623
rect 13863 15620 13875 15623
rect 13863 15592 15424 15620
rect 13863 15589 13875 15592
rect 13817 15583 13875 15589
rect 12084 15552 12112 15583
rect 12250 15552 12256 15564
rect 12084 15524 12256 15552
rect 12250 15512 12256 15524
rect 12308 15552 12314 15564
rect 12308 15524 12940 15552
rect 12308 15512 12314 15524
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 9824 15456 10701 15484
rect 9824 15444 9830 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 11698 15444 11704 15496
rect 11756 15484 11762 15496
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 11756 15456 12357 15484
rect 11756 15444 11762 15456
rect 12345 15453 12357 15456
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 12710 15444 12716 15496
rect 12768 15444 12774 15496
rect 12912 15493 12940 15524
rect 14734 15512 14740 15564
rect 14792 15552 14798 15564
rect 15197 15555 15255 15561
rect 15197 15552 15209 15555
rect 14792 15524 15209 15552
rect 14792 15512 14798 15524
rect 15197 15521 15209 15524
rect 15243 15521 15255 15555
rect 15197 15515 15255 15521
rect 15396 15496 15424 15592
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 13630 15444 13636 15496
rect 13688 15484 13694 15496
rect 14185 15487 14243 15493
rect 14185 15484 14197 15487
rect 13688 15456 14197 15484
rect 13688 15444 13694 15456
rect 14185 15453 14197 15456
rect 14231 15453 14243 15487
rect 14185 15447 14243 15453
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 10962 15425 10968 15428
rect 10956 15416 10968 15425
rect 10923 15388 10968 15416
rect 10956 15379 10968 15388
rect 10962 15376 10968 15379
rect 11020 15376 11026 15428
rect 13449 15419 13507 15425
rect 13449 15385 13461 15419
rect 13495 15416 13507 15419
rect 13814 15416 13820 15428
rect 13495 15388 13820 15416
rect 13495 15385 13507 15388
rect 13449 15379 13507 15385
rect 13814 15376 13820 15388
rect 13872 15376 13878 15428
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 13649 15351 13707 15357
rect 13649 15348 13661 15351
rect 12575 15320 13661 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 13649 15317 13661 15320
rect 13695 15348 13707 15351
rect 13906 15348 13912 15360
rect 13695 15320 13912 15348
rect 13695 15317 13707 15320
rect 13649 15311 13707 15317
rect 13906 15308 13912 15320
rect 13964 15348 13970 15360
rect 14660 15348 14688 15447
rect 15378 15444 15384 15496
rect 15436 15444 15442 15496
rect 15746 15444 15752 15496
rect 15804 15444 15810 15496
rect 15654 15376 15660 15428
rect 15712 15376 15718 15428
rect 13964 15320 14688 15348
rect 13964 15308 13970 15320
rect 1104 15258 28888 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 28888 15258
rect 1104 15184 28888 15206
rect 10962 15104 10968 15156
rect 11020 15144 11026 15156
rect 11609 15147 11667 15153
rect 11609 15144 11621 15147
rect 11020 15116 11621 15144
rect 11020 15104 11026 15116
rect 11609 15113 11621 15116
rect 11655 15113 11667 15147
rect 11609 15107 11667 15113
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 14277 15147 14335 15153
rect 14277 15144 14289 15147
rect 13872 15116 14289 15144
rect 13872 15104 13878 15116
rect 14277 15113 14289 15116
rect 14323 15144 14335 15147
rect 15286 15144 15292 15156
rect 14323 15116 15292 15144
rect 14323 15113 14335 15116
rect 14277 15107 14335 15113
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 9309 15011 9367 15017
rect 9309 14977 9321 15011
rect 9355 15008 9367 15011
rect 9766 15008 9772 15020
rect 9355 14980 9772 15008
rect 9355 14977 9367 14980
rect 9309 14971 9367 14977
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11664 14980 11805 15008
rect 11664 14968 11670 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 11882 14968 11888 15020
rect 11940 14968 11946 15020
rect 14826 14968 14832 15020
rect 14884 15008 14890 15020
rect 15105 15011 15163 15017
rect 15105 15008 15117 15011
rect 14884 14980 15117 15008
rect 14884 14968 14890 14980
rect 15105 14977 15117 14980
rect 15151 15008 15163 15011
rect 16574 15008 16580 15020
rect 15151 14980 16580 15008
rect 15151 14977 15163 14980
rect 15105 14971 15163 14977
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 23753 15011 23811 15017
rect 23753 14977 23765 15011
rect 23799 15008 23811 15011
rect 25130 15008 25136 15020
rect 23799 14980 25136 15008
rect 23799 14977 23811 14980
rect 23753 14971 23811 14977
rect 25130 14968 25136 14980
rect 25188 14968 25194 15020
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 11624 14940 11652 14968
rect 9732 14912 11652 14940
rect 13633 14943 13691 14949
rect 9732 14900 9738 14912
rect 13633 14909 13645 14943
rect 13679 14909 13691 14943
rect 13633 14903 13691 14909
rect 13648 14872 13676 14903
rect 14366 14900 14372 14952
rect 14424 14900 14430 14952
rect 14458 14900 14464 14952
rect 14516 14900 14522 14952
rect 14918 14900 14924 14952
rect 14976 14900 14982 14952
rect 24673 14943 24731 14949
rect 24673 14909 24685 14943
rect 24719 14940 24731 14943
rect 25406 14940 25412 14952
rect 24719 14912 25412 14940
rect 24719 14909 24731 14912
rect 24673 14903 24731 14909
rect 25406 14900 25412 14912
rect 25464 14900 25470 14952
rect 13909 14875 13967 14881
rect 13909 14872 13921 14875
rect 13648 14844 13921 14872
rect 13909 14841 13921 14844
rect 13955 14841 13967 14875
rect 13909 14835 13967 14841
rect 12986 14764 12992 14816
rect 13044 14764 13050 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15562 14804 15568 14816
rect 15335 14776 15568 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 23658 14764 23664 14816
rect 23716 14764 23722 14816
rect 24026 14764 24032 14816
rect 24084 14764 24090 14816
rect 1104 14714 28888 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 28888 14714
rect 1104 14640 28888 14662
rect 8478 14560 8484 14612
rect 8536 14560 8542 14612
rect 9766 14560 9772 14612
rect 9824 14560 9830 14612
rect 11330 14560 11336 14612
rect 11388 14560 11394 14612
rect 11882 14560 11888 14612
rect 11940 14600 11946 14612
rect 11977 14603 12035 14609
rect 11977 14600 11989 14603
rect 11940 14572 11989 14600
rect 11940 14560 11946 14572
rect 11977 14569 11989 14572
rect 12023 14569 12035 14603
rect 11977 14563 12035 14569
rect 13541 14603 13599 14609
rect 13541 14569 13553 14603
rect 13587 14600 13599 14603
rect 14366 14600 14372 14612
rect 13587 14572 14372 14600
rect 13587 14569 13599 14572
rect 13541 14563 13599 14569
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14976 14572 15117 14600
rect 14976 14560 14982 14572
rect 15105 14569 15117 14572
rect 15151 14569 15163 14603
rect 15105 14563 15163 14569
rect 25130 14560 25136 14612
rect 25188 14560 25194 14612
rect 25406 14560 25412 14612
rect 25464 14560 25470 14612
rect 8665 14535 8723 14541
rect 8665 14501 8677 14535
rect 8711 14532 8723 14535
rect 12526 14532 12532 14544
rect 8711 14504 12532 14532
rect 8711 14501 8723 14504
rect 8665 14495 8723 14501
rect 12526 14492 12532 14504
rect 12584 14492 12590 14544
rect 24121 14535 24179 14541
rect 24121 14501 24133 14535
rect 24167 14532 24179 14535
rect 24167 14504 24532 14532
rect 24167 14501 24179 14504
rect 24121 14495 24179 14501
rect 7098 14424 7104 14476
rect 7156 14464 7162 14476
rect 12621 14467 12679 14473
rect 7156 14436 8524 14464
rect 7156 14424 7162 14436
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14365 7803 14399
rect 7745 14359 7803 14365
rect 7374 14288 7380 14340
rect 7432 14328 7438 14340
rect 7760 14328 7788 14359
rect 7926 14356 7932 14408
rect 7984 14356 7990 14408
rect 8386 14356 8392 14408
rect 8444 14356 8450 14408
rect 8496 14405 8524 14436
rect 12621 14433 12633 14467
rect 12667 14464 12679 14467
rect 12710 14464 12716 14476
rect 12667 14436 12716 14464
rect 12667 14433 12679 14436
rect 12621 14427 12679 14433
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 24504 14473 24532 14504
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14464 13415 14467
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 13403 14436 15485 14464
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 15473 14433 15485 14436
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 20717 14467 20775 14473
rect 20717 14433 20729 14467
rect 20763 14464 20775 14467
rect 22741 14467 22799 14473
rect 22741 14464 22753 14467
rect 20763 14436 22753 14464
rect 20763 14433 20775 14436
rect 20717 14427 20775 14433
rect 22741 14433 22753 14436
rect 22787 14433 22799 14467
rect 22741 14427 22799 14433
rect 24489 14467 24547 14473
rect 24489 14433 24501 14467
rect 24535 14433 24547 14467
rect 25148 14464 25176 14560
rect 25148 14436 25636 14464
rect 24489 14427 24547 14433
rect 8481 14399 8539 14405
rect 8481 14365 8493 14399
rect 8527 14365 8539 14399
rect 8481 14359 8539 14365
rect 11057 14399 11115 14405
rect 11057 14365 11069 14399
rect 11103 14396 11115 14399
rect 11330 14396 11336 14408
rect 11103 14368 11336 14396
rect 11103 14365 11115 14368
rect 11057 14359 11115 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14396 13323 14399
rect 14274 14396 14280 14408
rect 13311 14368 14280 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 14424 14368 14473 14396
rect 14424 14356 14430 14368
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 15378 14356 15384 14408
rect 15436 14356 15442 14408
rect 15562 14356 15568 14408
rect 15620 14356 15626 14408
rect 19610 14356 19616 14408
rect 19668 14396 19674 14408
rect 20162 14396 20168 14408
rect 19668 14368 20168 14396
rect 19668 14356 19674 14368
rect 20162 14356 20168 14368
rect 20220 14396 20226 14408
rect 20732 14396 20760 14427
rect 20220 14368 20760 14396
rect 20993 14399 21051 14405
rect 20220 14356 20226 14368
rect 20993 14365 21005 14399
rect 21039 14365 21051 14399
rect 22756 14396 22784 14427
rect 24118 14396 24124 14408
rect 22756 14368 24124 14396
rect 20993 14359 21051 14365
rect 7432 14300 7788 14328
rect 7432 14288 7438 14300
rect 7558 14220 7564 14272
rect 7616 14220 7622 14272
rect 7760 14260 7788 14300
rect 8205 14331 8263 14337
rect 8205 14297 8217 14331
rect 8251 14328 8263 14331
rect 8294 14328 8300 14340
rect 8251 14300 8300 14328
rect 8251 14297 8263 14300
rect 8205 14291 8263 14297
rect 8294 14288 8300 14300
rect 8352 14288 8358 14340
rect 20254 14288 20260 14340
rect 20312 14328 20318 14340
rect 20450 14331 20508 14337
rect 20450 14328 20462 14331
rect 20312 14300 20462 14328
rect 20312 14288 20318 14300
rect 20450 14297 20462 14300
rect 20496 14297 20508 14331
rect 20450 14291 20508 14297
rect 9674 14260 9680 14272
rect 7760 14232 9680 14260
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 19337 14263 19395 14269
rect 19337 14229 19349 14263
rect 19383 14260 19395 14263
rect 20622 14260 20628 14272
rect 19383 14232 20628 14260
rect 19383 14229 19395 14232
rect 19337 14223 19395 14229
rect 20622 14220 20628 14232
rect 20680 14260 20686 14272
rect 21008 14260 21036 14359
rect 24118 14356 24124 14368
rect 24176 14356 24182 14408
rect 24854 14356 24860 14408
rect 24912 14396 24918 14408
rect 25608 14405 25636 14436
rect 25409 14399 25467 14405
rect 25409 14396 25421 14399
rect 24912 14368 25421 14396
rect 24912 14356 24918 14368
rect 25409 14365 25421 14368
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 25593 14399 25651 14405
rect 25593 14365 25605 14399
rect 25639 14365 25651 14399
rect 25593 14359 25651 14365
rect 28442 14356 28448 14408
rect 28500 14356 28506 14408
rect 23008 14331 23066 14337
rect 23008 14297 23020 14331
rect 23054 14328 23066 14331
rect 23198 14328 23204 14340
rect 23054 14300 23204 14328
rect 23054 14297 23066 14300
rect 23008 14291 23066 14297
rect 23198 14288 23204 14300
rect 23256 14288 23262 14340
rect 20680 14232 21036 14260
rect 20680 14220 20686 14232
rect 21634 14220 21640 14272
rect 21692 14220 21698 14272
rect 1104 14170 28888 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 28888 14170
rect 1104 14096 28888 14118
rect 7926 14016 7932 14068
rect 7984 14056 7990 14068
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 7984 14028 8769 14056
rect 7984 14016 7990 14028
rect 8757 14025 8769 14028
rect 8803 14056 8815 14059
rect 8803 14028 9904 14056
rect 8803 14025 8815 14028
rect 8757 14019 8815 14025
rect 9876 13997 9904 14028
rect 14366 14016 14372 14068
rect 14424 14016 14430 14068
rect 14737 14059 14795 14065
rect 14737 14025 14749 14059
rect 14783 14056 14795 14059
rect 15286 14056 15292 14068
rect 14783 14028 15292 14056
rect 14783 14025 14795 14028
rect 14737 14019 14795 14025
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 20254 14016 20260 14068
rect 20312 14016 20318 14068
rect 23198 14016 23204 14068
rect 23256 14016 23262 14068
rect 9861 13991 9919 13997
rect 9861 13957 9873 13991
rect 9907 13957 9919 13991
rect 9861 13951 9919 13957
rect 9953 13991 10011 13997
rect 9953 13957 9965 13991
rect 9999 13988 10011 13991
rect 10505 13991 10563 13997
rect 10505 13988 10517 13991
rect 9999 13960 10517 13988
rect 9999 13957 10011 13960
rect 9953 13951 10011 13957
rect 10505 13957 10517 13960
rect 10551 13957 10563 13991
rect 20438 13988 20444 14000
rect 10505 13951 10563 13957
rect 18984 13960 20444 13988
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7469 13855 7527 13861
rect 7469 13852 7481 13855
rect 7156 13824 7481 13852
rect 7156 13812 7162 13824
rect 7469 13821 7481 13824
rect 7515 13821 7527 13855
rect 7469 13815 7527 13821
rect 8110 13812 8116 13864
rect 8168 13812 8174 13864
rect 9784 13852 9812 13883
rect 10134 13880 10140 13932
rect 10192 13920 10198 13932
rect 10192 13892 10548 13920
rect 10192 13880 10198 13892
rect 10318 13852 10324 13864
rect 9784 13824 10324 13852
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10520 13852 10548 13892
rect 10594 13880 10600 13932
rect 10652 13920 10658 13932
rect 12434 13920 12440 13932
rect 10652 13892 12440 13920
rect 10652 13880 10658 13892
rect 12434 13880 12440 13892
rect 12492 13920 12498 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12492 13892 13001 13920
rect 12492 13880 12498 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 13256 13923 13314 13929
rect 13256 13889 13268 13923
rect 13302 13920 13314 13923
rect 13538 13920 13544 13932
rect 13302 13892 13544 13920
rect 13302 13889 13314 13892
rect 13256 13883 13314 13889
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 14918 13920 14924 13932
rect 14875 13892 14924 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 18984 13929 19012 13960
rect 20438 13948 20444 13960
rect 20496 13988 20502 14000
rect 20625 13991 20683 13997
rect 20625 13988 20637 13991
rect 20496 13960 20637 13988
rect 20496 13948 20502 13960
rect 20625 13957 20637 13960
rect 20671 13957 20683 13991
rect 20625 13951 20683 13957
rect 18969 13923 19027 13929
rect 18969 13920 18981 13923
rect 17512 13892 18981 13920
rect 10962 13852 10968 13864
rect 10520 13824 10968 13852
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11195 13824 12434 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 12406 13784 12434 13824
rect 12894 13784 12900 13796
rect 12406 13756 12900 13784
rect 12894 13744 12900 13756
rect 12952 13744 12958 13796
rect 17402 13744 17408 13796
rect 17460 13784 17466 13796
rect 17512 13784 17540 13892
rect 18969 13889 18981 13892
rect 19015 13889 19027 13923
rect 18969 13883 19027 13889
rect 19153 13923 19211 13929
rect 19153 13889 19165 13923
rect 19199 13920 19211 13923
rect 19199 13892 20024 13920
rect 19199 13889 19211 13892
rect 19153 13883 19211 13889
rect 18877 13855 18935 13861
rect 18877 13821 18889 13855
rect 18923 13852 18935 13855
rect 19337 13855 19395 13861
rect 18923 13824 19288 13852
rect 18923 13821 18935 13824
rect 18877 13815 18935 13821
rect 17460 13756 17540 13784
rect 19260 13784 19288 13824
rect 19337 13821 19349 13855
rect 19383 13852 19395 13855
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19383 13824 19625 13852
rect 19383 13821 19395 13824
rect 19337 13815 19395 13821
rect 19613 13821 19625 13824
rect 19659 13821 19671 13855
rect 19996 13852 20024 13892
rect 20530 13880 20536 13932
rect 20588 13880 20594 13932
rect 20806 13880 20812 13932
rect 20864 13920 20870 13932
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 20864 13892 21097 13920
rect 20864 13880 20870 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 24489 13923 24547 13929
rect 24489 13889 24501 13923
rect 24535 13920 24547 13923
rect 24946 13920 24952 13932
rect 24535 13892 24952 13920
rect 24535 13889 24547 13892
rect 24489 13883 24547 13889
rect 24946 13880 24952 13892
rect 25004 13880 25010 13932
rect 19996 13824 20852 13852
rect 19613 13815 19671 13821
rect 19978 13784 19984 13796
rect 19260 13756 19984 13784
rect 17460 13744 17466 13756
rect 19978 13744 19984 13756
rect 20036 13744 20042 13796
rect 20824 13793 20852 13824
rect 23750 13812 23756 13864
rect 23808 13812 23814 13864
rect 24394 13812 24400 13864
rect 24452 13812 24458 13864
rect 20809 13787 20867 13793
rect 20809 13753 20821 13787
rect 20855 13753 20867 13787
rect 20809 13747 20867 13753
rect 6914 13676 6920 13728
rect 6972 13676 6978 13728
rect 9585 13719 9643 13725
rect 9585 13685 9597 13719
rect 9631 13716 9643 13719
rect 10226 13716 10232 13728
rect 9631 13688 10232 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 24210 13676 24216 13728
rect 24268 13676 24274 13728
rect 1104 13626 28888 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 28888 13626
rect 1104 13552 28888 13574
rect 8110 13472 8116 13524
rect 8168 13472 8174 13524
rect 9766 13472 9772 13524
rect 9824 13512 9830 13524
rect 9824 13484 10272 13512
rect 9824 13472 9830 13484
rect 10134 13336 10140 13388
rect 10192 13336 10198 13388
rect 10244 13376 10272 13484
rect 10318 13472 10324 13524
rect 10376 13472 10382 13524
rect 11977 13515 12035 13521
rect 11977 13481 11989 13515
rect 12023 13512 12035 13515
rect 12710 13512 12716 13524
rect 12023 13484 12716 13512
rect 12023 13481 12035 13484
rect 11977 13475 12035 13481
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 13538 13472 13544 13524
rect 13596 13472 13602 13524
rect 15654 13404 15660 13456
rect 15712 13444 15718 13456
rect 23569 13447 23627 13453
rect 15712 13416 17540 13444
rect 15712 13404 15718 13416
rect 10594 13376 10600 13388
rect 10244 13348 10600 13376
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 16574 13336 16580 13388
rect 16632 13336 16638 13388
rect 17218 13376 17224 13388
rect 16684 13348 17224 13376
rect 6733 13311 6791 13317
rect 6733 13277 6745 13311
rect 6779 13308 6791 13311
rect 7282 13308 7288 13320
rect 6779 13280 7288 13308
rect 6779 13277 6791 13280
rect 6733 13271 6791 13277
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9582 13308 9588 13320
rect 9263 13280 9588 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 9674 13268 9680 13320
rect 9732 13268 9738 13320
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13308 10103 13311
rect 11330 13308 11336 13320
rect 10091 13280 11336 13308
rect 10091 13277 10103 13280
rect 10045 13271 10103 13277
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 16684 13317 16712 13348
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 17512 13385 17540 13416
rect 23569 13413 23581 13447
rect 23615 13444 23627 13447
rect 24394 13444 24400 13456
rect 23615 13416 24400 13444
rect 23615 13413 23627 13416
rect 23569 13407 23627 13413
rect 24394 13404 24400 13416
rect 24452 13404 24458 13456
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13345 17555 13379
rect 20717 13379 20775 13385
rect 20717 13376 20729 13379
rect 17497 13339 17555 13345
rect 20088 13348 20729 13376
rect 20088 13320 20116 13348
rect 20717 13345 20729 13348
rect 20763 13345 20775 13379
rect 20717 13339 20775 13345
rect 21726 13336 21732 13388
rect 21784 13376 21790 13388
rect 23109 13379 23167 13385
rect 23109 13376 23121 13379
rect 21784 13348 23121 13376
rect 21784 13336 21790 13348
rect 23109 13345 23121 13348
rect 23155 13345 23167 13379
rect 23109 13339 23167 13345
rect 13541 13311 13599 13317
rect 13541 13308 13553 13311
rect 13044 13280 13553 13308
rect 13044 13268 13050 13280
rect 13541 13277 13553 13280
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13308 13783 13311
rect 16669 13311 16727 13317
rect 13771 13280 14320 13308
rect 13771 13277 13783 13280
rect 13725 13271 13783 13277
rect 7006 13249 7012 13252
rect 7000 13203 7012 13249
rect 7006 13200 7012 13203
rect 7064 13200 7070 13252
rect 10870 13249 10876 13252
rect 9401 13243 9459 13249
rect 9401 13209 9413 13243
rect 9447 13240 9459 13243
rect 9769 13243 9827 13249
rect 9769 13240 9781 13243
rect 9447 13212 9781 13240
rect 9447 13209 9459 13212
rect 9401 13203 9459 13209
rect 9769 13209 9781 13212
rect 9815 13240 9827 13243
rect 9815 13212 10180 13240
rect 9815 13209 9827 13212
rect 9769 13203 9827 13209
rect 10152 13184 10180 13212
rect 10864 13203 10876 13249
rect 10870 13200 10876 13203
rect 10928 13200 10934 13252
rect 9950 13132 9956 13184
rect 10008 13132 10014 13184
rect 10134 13132 10140 13184
rect 10192 13132 10198 13184
rect 14292 13181 14320 13280
rect 16669 13277 16681 13311
rect 16715 13277 16727 13311
rect 16669 13271 16727 13277
rect 16850 13268 16856 13320
rect 16908 13308 16914 13320
rect 17313 13311 17371 13317
rect 17313 13308 17325 13311
rect 16908 13280 17325 13308
rect 16908 13268 16914 13280
rect 17313 13277 17325 13280
rect 17359 13277 17371 13311
rect 17313 13271 17371 13277
rect 17405 13311 17463 13317
rect 17405 13277 17417 13311
rect 17451 13277 17463 13311
rect 17405 13271 17463 13277
rect 17420 13240 17448 13271
rect 17586 13268 17592 13320
rect 17644 13268 17650 13320
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 19484 13280 19901 13308
rect 19484 13268 19490 13280
rect 19889 13277 19901 13280
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 20070 13268 20076 13320
rect 20128 13268 20134 13320
rect 20257 13311 20315 13317
rect 20257 13277 20269 13311
rect 20303 13277 20315 13311
rect 20257 13271 20315 13277
rect 16316 13212 17448 13240
rect 19352 13212 19932 13240
rect 16316 13184 16344 13212
rect 19352 13184 19380 13212
rect 14277 13175 14335 13181
rect 14277 13141 14289 13175
rect 14323 13172 14335 13175
rect 15194 13172 15200 13184
rect 14323 13144 15200 13172
rect 14323 13141 14335 13144
rect 14277 13135 14335 13141
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 16298 13132 16304 13184
rect 16356 13132 16362 13184
rect 17129 13175 17187 13181
rect 17129 13141 17141 13175
rect 17175 13172 17187 13175
rect 19334 13172 19340 13184
rect 17175 13144 19340 13172
rect 17175 13141 17187 13144
rect 17129 13135 17187 13141
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 19702 13132 19708 13184
rect 19760 13132 19766 13184
rect 19904 13172 19932 13212
rect 19978 13200 19984 13252
rect 20036 13200 20042 13252
rect 20272 13240 20300 13271
rect 20622 13268 20628 13320
rect 20680 13268 20686 13320
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 20732 13280 20821 13308
rect 20732 13240 20760 13280
rect 20809 13277 20821 13280
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 20898 13268 20904 13320
rect 20956 13268 20962 13320
rect 23201 13311 23259 13317
rect 23201 13277 23213 13311
rect 23247 13308 23259 13311
rect 23658 13308 23664 13320
rect 23247 13280 23664 13308
rect 23247 13277 23259 13280
rect 23201 13271 23259 13277
rect 23658 13268 23664 13280
rect 23716 13268 23722 13320
rect 20272 13212 20760 13240
rect 20272 13172 20300 13212
rect 19904 13144 20300 13172
rect 21085 13175 21143 13181
rect 21085 13141 21097 13175
rect 21131 13172 21143 13175
rect 23014 13172 23020 13184
rect 21131 13144 23020 13172
rect 21131 13141 21143 13144
rect 21085 13135 21143 13141
rect 23014 13132 23020 13144
rect 23072 13132 23078 13184
rect 23658 13132 23664 13184
rect 23716 13172 23722 13184
rect 23845 13175 23903 13181
rect 23845 13172 23857 13175
rect 23716 13144 23857 13172
rect 23716 13132 23722 13144
rect 23845 13141 23857 13144
rect 23891 13172 23903 13175
rect 23934 13172 23940 13184
rect 23891 13144 23940 13172
rect 23891 13141 23903 13144
rect 23845 13135 23903 13141
rect 23934 13132 23940 13144
rect 23992 13132 23998 13184
rect 1104 13082 28888 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 28888 13082
rect 1104 13008 28888 13030
rect 7006 12928 7012 12980
rect 7064 12928 7070 12980
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 8444 12940 8677 12968
rect 8444 12928 8450 12940
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 8665 12931 8723 12937
rect 6914 12900 6920 12912
rect 6748 12872 6920 12900
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 6748 12841 6776 12872
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 7374 12900 7380 12912
rect 7208 12872 7380 12900
rect 5905 12835 5963 12841
rect 5905 12832 5917 12835
rect 5592 12804 5917 12832
rect 5592 12792 5598 12804
rect 5905 12801 5917 12804
rect 5951 12832 5963 12835
rect 6733 12835 6791 12841
rect 5951 12804 6684 12832
rect 5951 12801 5963 12804
rect 5905 12795 5963 12801
rect 6086 12724 6092 12776
rect 6144 12724 6150 12776
rect 6656 12764 6684 12804
rect 6733 12801 6745 12835
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 7208 12832 7236 12872
rect 7374 12860 7380 12872
rect 7432 12860 7438 12912
rect 7558 12909 7564 12912
rect 7552 12900 7564 12909
rect 7519 12872 7564 12900
rect 7552 12863 7564 12872
rect 7558 12860 7564 12863
rect 7616 12860 7622 12912
rect 6871 12804 7236 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 6840 12764 6868 12795
rect 7282 12792 7288 12844
rect 7340 12792 7346 12844
rect 8680 12832 8708 12931
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 9585 12971 9643 12977
rect 9585 12968 9597 12971
rect 9180 12940 9597 12968
rect 9180 12928 9186 12940
rect 9585 12937 9597 12940
rect 9631 12937 9643 12971
rect 9585 12931 9643 12937
rect 10870 12928 10876 12980
rect 10928 12928 10934 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 11388 12940 12434 12968
rect 11388 12928 11394 12940
rect 9950 12860 9956 12912
rect 10008 12900 10014 12912
rect 12253 12903 12311 12909
rect 12253 12900 12265 12903
rect 10008 12872 12265 12900
rect 10008 12860 10014 12872
rect 12253 12869 12265 12872
rect 12299 12869 12311 12903
rect 12406 12900 12434 12940
rect 12894 12928 12900 12980
rect 12952 12968 12958 12980
rect 12989 12971 13047 12977
rect 12989 12968 13001 12971
rect 12952 12940 13001 12968
rect 12952 12928 12958 12940
rect 12989 12937 13001 12940
rect 13035 12937 13047 12971
rect 12989 12931 13047 12937
rect 16393 12971 16451 12977
rect 16393 12937 16405 12971
rect 16439 12968 16451 12971
rect 17221 12971 17279 12977
rect 17221 12968 17233 12971
rect 16439 12940 17233 12968
rect 16439 12937 16451 12940
rect 16393 12931 16451 12937
rect 17221 12937 17233 12940
rect 17267 12937 17279 12971
rect 17221 12931 17279 12937
rect 19797 12971 19855 12977
rect 19797 12937 19809 12971
rect 19843 12968 19855 12971
rect 20530 12968 20536 12980
rect 19843 12940 20536 12968
rect 19843 12937 19855 12940
rect 19797 12931 19855 12937
rect 20530 12928 20536 12940
rect 20588 12928 20594 12980
rect 20622 12928 20628 12980
rect 20680 12968 20686 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 20680 12940 22385 12968
rect 20680 12928 20686 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 22373 12931 22431 12937
rect 23566 12928 23572 12980
rect 23624 12968 23630 12980
rect 24121 12971 24179 12977
rect 24121 12968 24133 12971
rect 23624 12940 24133 12968
rect 23624 12928 23630 12940
rect 24121 12937 24133 12940
rect 24167 12968 24179 12971
rect 24854 12968 24860 12980
rect 24167 12940 24860 12968
rect 24167 12937 24179 12940
rect 24121 12931 24179 12937
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 24946 12928 24952 12980
rect 25004 12928 25010 12980
rect 17865 12903 17923 12909
rect 17865 12900 17877 12903
rect 12406 12872 12848 12900
rect 12253 12863 12311 12869
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8680 12804 8953 12832
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 10226 12792 10232 12844
rect 10284 12792 10290 12844
rect 6656 12736 6868 12764
rect 11606 12724 11612 12776
rect 11664 12724 11670 12776
rect 5718 12588 5724 12640
rect 5776 12588 5782 12640
rect 12268 12628 12296 12863
rect 12526 12792 12532 12844
rect 12584 12792 12590 12844
rect 12820 12841 12848 12872
rect 16040 12872 17877 12900
rect 12805 12835 12863 12841
rect 12805 12801 12817 12835
rect 12851 12801 12863 12835
rect 12805 12795 12863 12801
rect 15654 12792 15660 12844
rect 15712 12832 15718 12844
rect 16040 12841 16068 12872
rect 17865 12869 17877 12872
rect 17911 12869 17923 12903
rect 17865 12863 17923 12869
rect 19978 12860 19984 12912
rect 20036 12900 20042 12912
rect 20036 12872 21680 12900
rect 20036 12860 20042 12872
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15712 12804 16037 12832
rect 15712 12792 15718 12804
rect 16025 12801 16037 12804
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 17126 12792 17132 12844
rect 17184 12792 17190 12844
rect 17773 12835 17831 12841
rect 17773 12832 17785 12835
rect 17236 12804 17785 12832
rect 12618 12724 12624 12776
rect 12676 12724 12682 12776
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16298 12764 16304 12776
rect 16163 12736 16304 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16298 12724 16304 12736
rect 16356 12764 16362 12776
rect 17236 12764 17264 12804
rect 17773 12801 17785 12804
rect 17819 12801 17831 12835
rect 17773 12795 17831 12801
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 18506 12792 18512 12844
rect 18564 12792 18570 12844
rect 20456 12841 20484 12872
rect 21652 12844 21680 12872
rect 23750 12860 23756 12912
rect 23808 12860 23814 12912
rect 24210 12860 24216 12912
rect 24268 12860 24274 12912
rect 19429 12835 19487 12841
rect 19429 12801 19441 12835
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 20441 12835 20499 12841
rect 20441 12801 20453 12835
rect 20487 12801 20499 12835
rect 20441 12795 20499 12801
rect 16356 12736 17264 12764
rect 16356 12724 16362 12736
rect 17402 12724 17408 12776
rect 17460 12724 17466 12776
rect 19334 12724 19340 12776
rect 19392 12724 19398 12776
rect 19444 12764 19472 12795
rect 21266 12792 21272 12844
rect 21324 12792 21330 12844
rect 21634 12792 21640 12844
rect 21692 12832 21698 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21692 12804 22017 12832
rect 21692 12792 21698 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 20070 12764 20076 12776
rect 19444 12736 20076 12764
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 20349 12767 20407 12773
rect 20349 12733 20361 12767
rect 20395 12764 20407 12767
rect 21177 12767 21235 12773
rect 21177 12764 21189 12767
rect 20395 12736 21189 12764
rect 20395 12733 20407 12736
rect 20349 12727 20407 12733
rect 21177 12733 21189 12736
rect 21223 12764 21235 12767
rect 21726 12764 21732 12776
rect 21223 12736 21732 12764
rect 21223 12733 21235 12736
rect 21177 12727 21235 12733
rect 16666 12656 16672 12708
rect 16724 12696 16730 12708
rect 16724 12668 16896 12696
rect 16724 12656 16730 12668
rect 12529 12631 12587 12637
rect 12529 12628 12541 12631
rect 12268 12600 12541 12628
rect 12529 12597 12541 12600
rect 12575 12597 12587 12631
rect 12529 12591 12587 12597
rect 16758 12588 16764 12640
rect 16816 12588 16822 12640
rect 16868 12628 16896 12668
rect 17218 12656 17224 12708
rect 17276 12696 17282 12708
rect 18601 12699 18659 12705
rect 18601 12696 18613 12699
rect 17276 12668 18613 12696
rect 17276 12656 17282 12668
rect 18601 12665 18613 12668
rect 18647 12665 18659 12699
rect 18601 12659 18659 12665
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 20364 12696 20392 12727
rect 21726 12724 21732 12736
rect 21784 12724 21790 12776
rect 21818 12724 21824 12776
rect 21876 12764 21882 12776
rect 21913 12767 21971 12773
rect 21913 12764 21925 12767
rect 21876 12736 21925 12764
rect 21876 12724 21882 12736
rect 21913 12733 21925 12736
rect 21959 12733 21971 12767
rect 21913 12727 21971 12733
rect 19484 12668 20392 12696
rect 19484 12656 19490 12668
rect 20898 12656 20904 12708
rect 20956 12656 20962 12708
rect 21744 12696 21772 12724
rect 22204 12696 22232 12795
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 23109 12835 23167 12841
rect 23109 12832 23121 12835
rect 22520 12804 23121 12832
rect 22520 12792 22526 12804
rect 23109 12801 23121 12804
rect 23155 12801 23167 12835
rect 23109 12795 23167 12801
rect 23658 12792 23664 12844
rect 23716 12832 23722 12844
rect 23845 12835 23903 12841
rect 23845 12832 23857 12835
rect 23716 12804 23857 12832
rect 23716 12792 23722 12804
rect 23845 12801 23857 12804
rect 23891 12801 23903 12835
rect 23845 12795 23903 12801
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12832 23995 12835
rect 24026 12832 24032 12844
rect 23983 12804 24032 12832
rect 23983 12801 23995 12804
rect 23937 12795 23995 12801
rect 24026 12792 24032 12804
rect 24084 12792 24090 12844
rect 24489 12835 24547 12841
rect 24489 12801 24501 12835
rect 24535 12801 24547 12835
rect 24489 12795 24547 12801
rect 23014 12724 23020 12776
rect 23072 12764 23078 12776
rect 23072 12736 23796 12764
rect 23072 12724 23078 12736
rect 21744 12668 22232 12696
rect 23474 12656 23480 12708
rect 23532 12656 23538 12708
rect 23768 12696 23796 12736
rect 24504 12696 24532 12795
rect 24578 12792 24584 12844
rect 24636 12792 24642 12844
rect 24762 12792 24768 12844
rect 24820 12792 24826 12844
rect 23768 12668 24532 12696
rect 17402 12628 17408 12640
rect 16868 12600 17408 12628
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 18230 12588 18236 12640
rect 18288 12588 18294 12640
rect 1104 12538 28888 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 28888 12538
rect 1104 12464 28888 12486
rect 9398 12424 9404 12436
rect 9140 12396 9404 12424
rect 8665 12359 8723 12365
rect 8665 12325 8677 12359
rect 8711 12356 8723 12359
rect 9140 12356 9168 12396
rect 9398 12384 9404 12396
rect 9456 12424 9462 12436
rect 9456 12396 10916 12424
rect 9456 12384 9462 12396
rect 8711 12328 9168 12356
rect 10888 12356 10916 12396
rect 11330 12384 11336 12436
rect 11388 12384 11394 12436
rect 11606 12384 11612 12436
rect 11664 12384 11670 12436
rect 12618 12424 12624 12436
rect 11716 12396 12624 12424
rect 11716 12356 11744 12396
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 14458 12384 14464 12436
rect 14516 12424 14522 12436
rect 16666 12424 16672 12436
rect 14516 12396 16672 12424
rect 14516 12384 14522 12396
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 16850 12384 16856 12436
rect 16908 12384 16914 12436
rect 18325 12427 18383 12433
rect 18325 12393 18337 12427
rect 18371 12424 18383 12427
rect 18506 12424 18512 12436
rect 18371 12396 18512 12424
rect 18371 12393 18383 12396
rect 18325 12387 18383 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 16868 12356 16896 12384
rect 10888 12328 11744 12356
rect 15764 12328 16896 12356
rect 8711 12325 8723 12328
rect 8665 12319 8723 12325
rect 9140 12297 9168 12328
rect 15764 12297 15792 12328
rect 18046 12316 18052 12368
rect 18104 12356 18110 12368
rect 18601 12359 18659 12365
rect 18601 12356 18613 12359
rect 18104 12328 18613 12356
rect 18104 12316 18110 12328
rect 18601 12325 18613 12328
rect 18647 12325 18659 12359
rect 23566 12356 23572 12368
rect 18601 12319 18659 12325
rect 23308 12328 23572 12356
rect 9125 12291 9183 12297
rect 9125 12257 9137 12291
rect 9171 12257 9183 12291
rect 9125 12251 9183 12257
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 16758 12248 16764 12300
rect 16816 12288 16822 12300
rect 16853 12291 16911 12297
rect 16853 12288 16865 12291
rect 16816 12260 16865 12288
rect 16816 12248 16822 12260
rect 16853 12257 16865 12260
rect 16899 12257 16911 12291
rect 18230 12288 18236 12300
rect 16853 12251 16911 12257
rect 17420 12260 18236 12288
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 5629 12223 5687 12229
rect 5629 12220 5641 12223
rect 5500 12192 5641 12220
rect 5500 12180 5506 12192
rect 5629 12189 5641 12192
rect 5675 12220 5687 12223
rect 7282 12220 7288 12232
rect 5675 12192 7288 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 7282 12180 7288 12192
rect 7340 12220 7346 12232
rect 7340 12192 8248 12220
rect 7340 12180 7346 12192
rect 5718 12112 5724 12164
rect 5776 12152 5782 12164
rect 5874 12155 5932 12161
rect 5874 12152 5886 12155
rect 5776 12124 5886 12152
rect 5776 12112 5782 12124
rect 5874 12121 5886 12124
rect 5920 12121 5932 12155
rect 5874 12115 5932 12121
rect 7552 12155 7610 12161
rect 7552 12121 7564 12155
rect 7598 12152 7610 12155
rect 7926 12152 7932 12164
rect 7598 12124 7932 12152
rect 7598 12121 7610 12124
rect 7552 12115 7610 12121
rect 7926 12112 7932 12124
rect 7984 12112 7990 12164
rect 8220 12152 8248 12192
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10594 12220 10600 12232
rect 10008 12192 10600 12220
rect 10008 12180 10014 12192
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 12492 12192 13001 12220
rect 12492 12180 12498 12192
rect 12989 12189 13001 12192
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 17420 12220 17448 12260
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 18340 12260 18981 12288
rect 15703 12192 17448 12220
rect 17773 12223 17831 12229
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 17773 12189 17785 12223
rect 17819 12220 17831 12223
rect 17954 12220 17960 12232
rect 17819 12192 17960 12220
rect 17819 12189 17831 12192
rect 17773 12183 17831 12189
rect 17954 12180 17960 12192
rect 18012 12220 18018 12232
rect 18340 12220 18368 12260
rect 18969 12257 18981 12260
rect 19015 12257 19027 12291
rect 18969 12251 19027 12257
rect 19702 12248 19708 12300
rect 19760 12248 19766 12300
rect 20438 12248 20444 12300
rect 20496 12288 20502 12300
rect 23308 12297 23336 12328
rect 23566 12316 23572 12328
rect 23624 12316 23630 12368
rect 23845 12359 23903 12365
rect 23845 12325 23857 12359
rect 23891 12356 23903 12359
rect 23891 12328 24532 12356
rect 23891 12325 23903 12328
rect 23845 12319 23903 12325
rect 20809 12291 20867 12297
rect 20809 12288 20821 12291
rect 20496 12260 20821 12288
rect 20496 12248 20502 12260
rect 20809 12257 20821 12260
rect 20855 12288 20867 12291
rect 23293 12291 23351 12297
rect 23293 12288 23305 12291
rect 20855 12260 23305 12288
rect 20855 12257 20867 12260
rect 20809 12251 20867 12257
rect 23293 12257 23305 12260
rect 23339 12257 23351 12291
rect 23293 12251 23351 12257
rect 23385 12291 23443 12297
rect 23385 12257 23397 12291
rect 23431 12288 23443 12291
rect 23474 12288 23480 12300
rect 23431 12260 23480 12288
rect 23431 12257 23443 12260
rect 23385 12251 23443 12257
rect 23474 12248 23480 12260
rect 23532 12248 23538 12300
rect 24504 12297 24532 12328
rect 24489 12291 24547 12297
rect 24489 12257 24501 12291
rect 24535 12257 24547 12291
rect 24489 12251 24547 12257
rect 18012 12192 18368 12220
rect 18785 12223 18843 12229
rect 18012 12180 18018 12192
rect 18785 12189 18797 12223
rect 18831 12220 18843 12223
rect 19426 12220 19432 12232
rect 18831 12192 19432 12220
rect 18831 12189 18843 12192
rect 18785 12183 18843 12189
rect 9968 12152 9996 12180
rect 10226 12161 10232 12164
rect 8220 12124 9996 12152
rect 10220 12115 10232 12161
rect 10226 12112 10232 12115
rect 10284 12112 10290 12164
rect 10686 12112 10692 12164
rect 10744 12152 10750 12164
rect 12722 12155 12780 12161
rect 12722 12152 12734 12155
rect 10744 12124 12734 12152
rect 10744 12112 10750 12124
rect 12722 12121 12734 12124
rect 12768 12121 12780 12155
rect 12722 12115 12780 12121
rect 17862 12112 17868 12164
rect 17920 12152 17926 12164
rect 18800 12152 18828 12183
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 19613 12223 19671 12229
rect 19613 12189 19625 12223
rect 19659 12220 19671 12223
rect 20898 12220 20904 12232
rect 19659 12192 20904 12220
rect 19659 12189 19671 12192
rect 19613 12183 19671 12189
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21818 12180 21824 12232
rect 21876 12180 21882 12232
rect 22738 12180 22744 12232
rect 22796 12180 22802 12232
rect 20717 12155 20775 12161
rect 20717 12152 20729 12155
rect 17920 12124 18828 12152
rect 19996 12124 20729 12152
rect 17920 12112 17926 12124
rect 7006 12044 7012 12096
rect 7064 12044 7070 12096
rect 9677 12087 9735 12093
rect 9677 12053 9689 12087
rect 9723 12084 9735 12087
rect 10042 12084 10048 12096
rect 9723 12056 10048 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 16022 12044 16028 12096
rect 16080 12044 16086 12096
rect 16298 12044 16304 12096
rect 16356 12044 16362 12096
rect 19996 12093 20024 12124
rect 20717 12121 20729 12124
rect 20763 12121 20775 12155
rect 20717 12115 20775 12121
rect 22278 12112 22284 12164
rect 22336 12152 22342 12164
rect 23477 12155 23535 12161
rect 23477 12152 23489 12155
rect 22336 12124 23489 12152
rect 22336 12112 22342 12124
rect 23477 12121 23489 12124
rect 23523 12121 23535 12155
rect 23477 12115 23535 12121
rect 19981 12087 20039 12093
rect 19981 12053 19993 12087
rect 20027 12053 20039 12087
rect 19981 12047 20039 12053
rect 20254 12044 20260 12096
rect 20312 12044 20318 12096
rect 20625 12087 20683 12093
rect 20625 12053 20637 12087
rect 20671 12084 20683 12087
rect 21174 12084 21180 12096
rect 20671 12056 21180 12084
rect 20671 12053 20683 12056
rect 20625 12047 20683 12053
rect 21174 12044 21180 12056
rect 21232 12044 21238 12096
rect 21269 12087 21327 12093
rect 21269 12053 21281 12087
rect 21315 12084 21327 12087
rect 21450 12084 21456 12096
rect 21315 12056 21456 12084
rect 21315 12053 21327 12056
rect 21269 12047 21327 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 22186 12044 22192 12096
rect 22244 12044 22250 12096
rect 25130 12044 25136 12096
rect 25188 12044 25194 12096
rect 1104 11994 28888 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 28888 11994
rect 1104 11920 28888 11942
rect 6086 11840 6092 11892
rect 6144 11880 6150 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 6144 11852 6469 11880
rect 6144 11840 6150 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 8352 11852 8585 11880
rect 8352 11840 8358 11852
rect 8573 11849 8585 11852
rect 8619 11849 8631 11883
rect 8573 11843 8631 11849
rect 16761 11883 16819 11889
rect 16761 11849 16773 11883
rect 16807 11880 16819 11883
rect 16850 11880 16856 11892
rect 16807 11852 16856 11880
rect 16807 11849 16819 11852
rect 16761 11843 16819 11849
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 17586 11840 17592 11892
rect 17644 11840 17650 11892
rect 20993 11883 21051 11889
rect 20993 11849 21005 11883
rect 21039 11880 21051 11883
rect 21818 11880 21824 11892
rect 21039 11852 21824 11880
rect 21039 11849 21051 11852
rect 20993 11843 21051 11849
rect 21818 11840 21824 11852
rect 21876 11840 21882 11892
rect 22462 11840 22468 11892
rect 22520 11840 22526 11892
rect 22738 11840 22744 11892
rect 22796 11840 22802 11892
rect 24762 11880 24768 11892
rect 23768 11852 24768 11880
rect 18138 11812 18144 11824
rect 17144 11784 18144 11812
rect 5534 11704 5540 11756
rect 5592 11704 5598 11756
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11744 5687 11747
rect 5902 11744 5908 11756
rect 5675 11716 5908 11744
rect 5675 11713 5687 11716
rect 5629 11707 5687 11713
rect 5902 11704 5908 11716
rect 5960 11704 5966 11756
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 9697 11747 9755 11753
rect 9697 11713 9709 11747
rect 9743 11744 9755 11747
rect 9858 11744 9864 11756
rect 9743 11716 9864 11744
rect 9743 11713 9755 11716
rect 9697 11707 9755 11713
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 9950 11704 9956 11756
rect 10008 11704 10014 11756
rect 11241 11747 11299 11753
rect 11241 11713 11253 11747
rect 11287 11744 11299 11747
rect 11330 11744 11336 11756
rect 11287 11716 11336 11744
rect 11287 11713 11299 11716
rect 11241 11707 11299 11713
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 14366 11704 14372 11756
rect 14424 11704 14430 11756
rect 14458 11704 14464 11756
rect 14516 11744 14522 11756
rect 14553 11747 14611 11753
rect 14553 11744 14565 11747
rect 14516 11716 14565 11744
rect 14516 11704 14522 11716
rect 14553 11713 14565 11716
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 15194 11704 15200 11756
rect 15252 11744 15258 11756
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 15252 11716 15669 11744
rect 15252 11704 15258 11716
rect 15657 11713 15669 11716
rect 15703 11713 15715 11747
rect 15657 11707 15715 11713
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16298 11744 16304 11756
rect 15887 11716 16304 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 7101 11679 7159 11685
rect 7101 11676 7113 11679
rect 6880 11648 7113 11676
rect 6880 11636 6886 11648
rect 7101 11645 7113 11648
rect 7147 11676 7159 11679
rect 8478 11676 8484 11688
rect 7147 11648 8484 11676
rect 7147 11645 7159 11648
rect 7101 11639 7159 11645
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 14332 11648 14657 11676
rect 14332 11636 14338 11648
rect 14645 11645 14657 11648
rect 14691 11676 14703 11679
rect 14918 11676 14924 11688
rect 14691 11648 14924 11676
rect 14691 11645 14703 11648
rect 14645 11639 14703 11645
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 15672 11676 15700 11707
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 17144 11753 17172 11784
rect 18138 11772 18144 11784
rect 18196 11772 18202 11824
rect 21266 11772 21272 11824
rect 21324 11812 21330 11824
rect 21361 11815 21419 11821
rect 21361 11812 21373 11815
rect 21324 11784 21373 11812
rect 21324 11772 21330 11784
rect 21361 11781 21373 11784
rect 21407 11781 21419 11815
rect 21361 11775 21419 11781
rect 22005 11815 22063 11821
rect 22005 11781 22017 11815
rect 22051 11812 22063 11815
rect 23768 11812 23796 11852
rect 24762 11840 24768 11852
rect 24820 11880 24826 11892
rect 24857 11883 24915 11889
rect 24857 11880 24869 11883
rect 24820 11852 24869 11880
rect 24820 11840 24826 11852
rect 24857 11849 24869 11852
rect 24903 11849 24915 11883
rect 24857 11843 24915 11849
rect 22051 11784 23796 11812
rect 23876 11815 23934 11821
rect 22051 11781 22063 11784
rect 22005 11775 22063 11781
rect 23876 11781 23888 11815
rect 23922 11812 23934 11815
rect 25225 11815 25283 11821
rect 25225 11812 25237 11815
rect 23922 11784 25237 11812
rect 23922 11781 23934 11784
rect 23876 11775 23934 11781
rect 25225 11781 25237 11784
rect 25271 11781 25283 11815
rect 25225 11775 25283 11781
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17773 11747 17831 11753
rect 17773 11713 17785 11747
rect 17819 11744 17831 11747
rect 17862 11744 17868 11756
rect 17819 11716 17868 11744
rect 17819 11713 17831 11716
rect 17773 11707 17831 11713
rect 16117 11679 16175 11685
rect 16117 11676 16129 11679
rect 15672 11648 16129 11676
rect 16117 11645 16129 11648
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 16132 11608 16160 11639
rect 16574 11636 16580 11688
rect 16632 11676 16638 11688
rect 17037 11679 17095 11685
rect 17037 11676 17049 11679
rect 16632 11648 17049 11676
rect 16632 11636 16638 11648
rect 17037 11645 17049 11648
rect 17083 11676 17095 11679
rect 17788 11676 17816 11707
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 19886 11753 19892 11756
rect 19880 11707 19892 11753
rect 19886 11704 19892 11707
rect 19944 11704 19950 11756
rect 21450 11704 21456 11756
rect 21508 11704 21514 11756
rect 21726 11704 21732 11756
rect 21784 11744 21790 11756
rect 21784 11716 24072 11744
rect 21784 11704 21790 11716
rect 17083 11648 17816 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 18046 11636 18052 11688
rect 18104 11636 18110 11688
rect 19610 11636 19616 11688
rect 19668 11636 19674 11688
rect 24044 11676 24072 11716
rect 24118 11704 24124 11756
rect 24176 11704 24182 11756
rect 24673 11747 24731 11753
rect 24673 11744 24685 11747
rect 24228 11716 24685 11744
rect 24228 11676 24256 11716
rect 24673 11713 24685 11716
rect 24719 11713 24731 11747
rect 24673 11707 24731 11713
rect 25130 11704 25136 11756
rect 25188 11704 25194 11756
rect 25317 11747 25375 11753
rect 25317 11713 25329 11747
rect 25363 11744 25375 11747
rect 25593 11747 25651 11753
rect 25593 11744 25605 11747
rect 25363 11716 25605 11744
rect 25363 11713 25375 11716
rect 25317 11707 25375 11713
rect 25593 11713 25605 11716
rect 25639 11713 25651 11747
rect 25593 11707 25651 11713
rect 24044 11648 24256 11676
rect 24486 11636 24492 11688
rect 24544 11636 24550 11688
rect 24762 11636 24768 11688
rect 24820 11676 24826 11688
rect 25332 11676 25360 11707
rect 24820 11648 25360 11676
rect 24820 11636 24826 11648
rect 19518 11608 19524 11620
rect 16132 11580 19524 11608
rect 19518 11568 19524 11580
rect 19576 11568 19582 11620
rect 22373 11611 22431 11617
rect 22373 11577 22385 11611
rect 22419 11577 22431 11611
rect 22373 11571 22431 11577
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 5776 11512 5825 11540
rect 5776 11500 5782 11512
rect 5813 11509 5825 11512
rect 5859 11509 5871 11543
rect 5813 11503 5871 11509
rect 7653 11543 7711 11549
rect 7653 11509 7665 11543
rect 7699 11540 7711 11543
rect 8294 11540 8300 11552
rect 7699 11512 8300 11540
rect 7699 11509 7711 11512
rect 7653 11503 7711 11509
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 10594 11500 10600 11552
rect 10652 11500 10658 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 14148 11512 14197 11540
rect 14148 11500 14154 11512
rect 14185 11509 14197 11512
rect 14231 11509 14243 11543
rect 14185 11503 14243 11509
rect 15838 11500 15844 11552
rect 15896 11500 15902 11552
rect 17954 11500 17960 11552
rect 18012 11500 18018 11552
rect 19536 11540 19564 11568
rect 20806 11540 20812 11552
rect 19536 11512 20812 11540
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 22094 11500 22100 11552
rect 22152 11540 22158 11552
rect 22388 11540 22416 11571
rect 24578 11540 24584 11552
rect 22152 11512 24584 11540
rect 22152 11500 22158 11512
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 1104 11450 28888 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 28888 11450
rect 1104 11376 28888 11398
rect 6822 11296 6828 11348
rect 6880 11296 6886 11348
rect 7926 11296 7932 11348
rect 7984 11296 7990 11348
rect 9585 11339 9643 11345
rect 9585 11305 9597 11339
rect 9631 11336 9643 11339
rect 9674 11336 9680 11348
rect 9631 11308 9680 11336
rect 9631 11305 9643 11308
rect 9585 11299 9643 11305
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10597 11339 10655 11345
rect 10597 11305 10609 11339
rect 10643 11336 10655 11339
rect 10686 11336 10692 11348
rect 10643 11308 10692 11336
rect 10643 11305 10655 11308
rect 10597 11299 10655 11305
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 14918 11296 14924 11348
rect 14976 11296 14982 11348
rect 16022 11296 16028 11348
rect 16080 11336 16086 11348
rect 16761 11339 16819 11345
rect 16080 11308 16574 11336
rect 16080 11296 16086 11308
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 9033 11271 9091 11277
rect 9033 11268 9045 11271
rect 7064 11240 9045 11268
rect 7064 11228 7070 11240
rect 9033 11237 9045 11240
rect 9079 11237 9091 11271
rect 9033 11231 9091 11237
rect 13817 11271 13875 11277
rect 13817 11237 13829 11271
rect 13863 11268 13875 11271
rect 13863 11240 14320 11268
rect 13863 11237 13875 11240
rect 13817 11231 13875 11237
rect 5442 11160 5448 11212
rect 5500 11160 5506 11212
rect 8294 11160 8300 11212
rect 8352 11160 8358 11212
rect 10042 11160 10048 11212
rect 10100 11200 10106 11212
rect 10229 11203 10287 11209
rect 10229 11200 10241 11203
rect 10100 11172 10241 11200
rect 10100 11160 10106 11172
rect 10229 11169 10241 11172
rect 10275 11169 10287 11203
rect 10229 11163 10287 11169
rect 12434 11160 12440 11212
rect 12492 11160 12498 11212
rect 14292 11209 14320 11240
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11169 14335 11203
rect 16546 11200 16574 11308
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 17954 11336 17960 11348
rect 16807 11308 17960 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 17954 11296 17960 11308
rect 18012 11296 18018 11348
rect 18138 11296 18144 11348
rect 18196 11296 18202 11348
rect 19886 11296 19892 11348
rect 19944 11296 19950 11348
rect 22094 11296 22100 11348
rect 22152 11296 22158 11348
rect 22278 11296 22284 11348
rect 22336 11336 22342 11348
rect 22465 11339 22523 11345
rect 22465 11336 22477 11339
rect 22336 11308 22477 11336
rect 22336 11296 22342 11308
rect 22465 11305 22477 11308
rect 22511 11305 22523 11339
rect 22465 11299 22523 11305
rect 23842 11296 23848 11348
rect 23900 11296 23906 11348
rect 17402 11228 17408 11280
rect 17460 11268 17466 11280
rect 17460 11240 17632 11268
rect 17460 11228 17466 11240
rect 17604 11209 17632 11240
rect 20806 11228 20812 11280
rect 20864 11268 20870 11280
rect 23477 11271 23535 11277
rect 23477 11268 23489 11271
rect 20864 11240 23489 11268
rect 20864 11228 20870 11240
rect 23477 11237 23489 11240
rect 23523 11268 23535 11271
rect 23658 11268 23664 11280
rect 23523 11240 23664 11268
rect 23523 11237 23535 11240
rect 23477 11231 23535 11237
rect 23658 11228 23664 11240
rect 23716 11268 23722 11280
rect 24489 11271 24547 11277
rect 24489 11268 24501 11271
rect 23716 11240 24501 11268
rect 23716 11228 23722 11240
rect 24489 11237 24501 11240
rect 24535 11268 24547 11271
rect 24762 11268 24768 11280
rect 24535 11240 24768 11268
rect 24535 11237 24547 11240
rect 24489 11231 24547 11237
rect 24762 11228 24768 11240
rect 24820 11228 24826 11280
rect 17497 11203 17555 11209
rect 17497 11200 17509 11203
rect 16546 11172 17509 11200
rect 14277 11163 14335 11169
rect 17497 11169 17509 11172
rect 17543 11169 17555 11203
rect 17497 11163 17555 11169
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11169 17647 11203
rect 19610 11200 19616 11212
rect 17589 11163 17647 11169
rect 18156 11172 19616 11200
rect 5718 11141 5724 11144
rect 5712 11132 5724 11141
rect 5679 11104 5724 11132
rect 5712 11095 5724 11104
rect 5718 11092 5724 11095
rect 5776 11092 5782 11144
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 7432 11104 8125 11132
rect 7432 11092 7438 11104
rect 8113 11101 8125 11104
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 8444 11104 9321 11132
rect 8444 11092 8450 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 9640 11104 10425 11132
rect 9640 11092 9646 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 16206 11132 16212 11144
rect 15427 11104 16212 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 16206 11092 16212 11104
rect 16264 11132 16270 11144
rect 18156 11132 18184 11172
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 20717 11203 20775 11209
rect 20717 11200 20729 11203
rect 20312 11172 20729 11200
rect 20312 11160 20318 11172
rect 20717 11169 20729 11172
rect 20763 11169 20775 11203
rect 20717 11163 20775 11169
rect 16264 11104 18184 11132
rect 16264 11092 16270 11104
rect 18230 11092 18236 11144
rect 18288 11092 18294 11144
rect 19518 11092 19524 11144
rect 19576 11132 19582 11144
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 19576 11104 19717 11132
rect 19576 11092 19582 11104
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 19889 11135 19947 11141
rect 19889 11101 19901 11135
rect 19935 11132 19947 11135
rect 20165 11135 20223 11141
rect 20165 11132 20177 11135
rect 19935 11104 20177 11132
rect 19935 11101 19947 11104
rect 19889 11095 19947 11101
rect 20165 11101 20177 11104
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 21726 11092 21732 11144
rect 21784 11092 21790 11144
rect 21913 11135 21971 11141
rect 21913 11101 21925 11135
rect 21959 11132 21971 11135
rect 22186 11132 22192 11144
rect 21959 11104 22192 11132
rect 21959 11101 21971 11104
rect 21913 11095 21971 11101
rect 22186 11092 22192 11104
rect 22244 11132 22250 11144
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 22244 11104 22569 11132
rect 22244 11092 22250 11104
rect 22557 11101 22569 11104
rect 22603 11132 22615 11135
rect 24486 11132 24492 11144
rect 22603 11104 24492 11132
rect 22603 11101 22615 11104
rect 22557 11095 22615 11101
rect 24486 11092 24492 11104
rect 24544 11092 24550 11144
rect 8478 11024 8484 11076
rect 8536 11064 8542 11076
rect 9217 11067 9275 11073
rect 9217 11064 9229 11067
rect 8536 11036 9229 11064
rect 8536 11024 8542 11036
rect 9217 11033 9229 11036
rect 9263 11033 9275 11067
rect 9217 11027 9275 11033
rect 12704 11067 12762 11073
rect 12704 11033 12716 11067
rect 12750 11064 12762 11067
rect 13446 11064 13452 11076
rect 12750 11036 13452 11064
rect 12750 11033 12762 11036
rect 12704 11027 12762 11033
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 15648 11067 15706 11073
rect 15648 11033 15660 11067
rect 15694 11064 15706 11067
rect 15838 11064 15844 11076
rect 15694 11036 15844 11064
rect 15694 11033 15706 11036
rect 15648 11027 15706 11033
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 17405 11067 17463 11073
rect 17405 11033 17417 11067
rect 17451 11064 17463 11067
rect 18138 11064 18144 11076
rect 17451 11036 18144 11064
rect 17451 11033 17463 11036
rect 17405 11027 17463 11033
rect 18138 11024 18144 11036
rect 18196 11024 18202 11076
rect 23201 11067 23259 11073
rect 23201 11033 23213 11067
rect 23247 11064 23259 11067
rect 23842 11064 23848 11076
rect 23247 11036 23848 11064
rect 23247 11033 23259 11036
rect 23201 11027 23259 11033
rect 23842 11024 23848 11036
rect 23900 11064 23906 11076
rect 28258 11064 28264 11076
rect 23900 11036 28264 11064
rect 23900 11024 23906 11036
rect 28258 11024 28264 11036
rect 28316 11024 28322 11076
rect 17034 10956 17040 11008
rect 17092 10956 17098 11008
rect 1104 10906 28888 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 28888 10906
rect 1104 10832 28888 10854
rect 9493 10795 9551 10801
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 9858 10792 9864 10804
rect 9539 10764 9864 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 13446 10752 13452 10804
rect 13504 10752 13510 10804
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 14918 10792 14924 10804
rect 14599 10764 14924 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 18509 10795 18567 10801
rect 18509 10792 18521 10795
rect 18288 10764 18521 10792
rect 18288 10752 18294 10764
rect 18509 10761 18521 10764
rect 18555 10761 18567 10795
rect 18509 10755 18567 10761
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 19981 10795 20039 10801
rect 19981 10792 19993 10795
rect 19576 10764 19993 10792
rect 19576 10752 19582 10764
rect 19981 10761 19993 10764
rect 20027 10761 20039 10795
rect 19981 10755 20039 10761
rect 14369 10727 14427 10733
rect 14369 10693 14381 10727
rect 14415 10724 14427 10727
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 14415 10696 15025 10724
rect 14415 10693 14427 10696
rect 14369 10687 14427 10693
rect 15013 10693 15025 10696
rect 15059 10724 15071 10727
rect 15194 10724 15200 10736
rect 15059 10696 15200 10724
rect 15059 10693 15071 10696
rect 15013 10687 15071 10693
rect 15194 10684 15200 10696
rect 15252 10684 15258 10736
rect 9674 10616 9680 10668
rect 9732 10616 9738 10668
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10656 9919 10659
rect 10594 10656 10600 10668
rect 9907 10628 10600 10656
rect 9907 10625 9919 10628
rect 9861 10619 9919 10625
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 14090 10616 14096 10668
rect 14148 10616 14154 10668
rect 14458 10616 14464 10668
rect 14516 10656 14522 10668
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14516 10628 14657 10656
rect 14516 10616 14522 10628
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 17034 10616 17040 10668
rect 17092 10656 17098 10668
rect 17313 10659 17371 10665
rect 17313 10656 17325 10659
rect 17092 10628 17325 10656
rect 17092 10616 17098 10628
rect 17313 10625 17325 10628
rect 17359 10625 17371 10659
rect 17313 10619 17371 10625
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10656 17923 10659
rect 18046 10656 18052 10668
rect 17911 10628 18052 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 14366 10480 14372 10532
rect 14424 10480 14430 10532
rect 15930 10412 15936 10464
rect 15988 10452 15994 10464
rect 16761 10455 16819 10461
rect 16761 10452 16773 10455
rect 15988 10424 16773 10452
rect 15988 10412 15994 10424
rect 16761 10421 16773 10424
rect 16807 10421 16819 10455
rect 16761 10415 16819 10421
rect 1104 10362 28888 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 28888 10362
rect 1104 10288 28888 10310
rect 17589 10251 17647 10257
rect 17589 10217 17601 10251
rect 17635 10248 17647 10251
rect 18046 10248 18052 10260
rect 17635 10220 18052 10248
rect 17635 10217 17647 10220
rect 17589 10211 17647 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 16206 10072 16212 10124
rect 16264 10072 16270 10124
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15746 10044 15752 10056
rect 15252 10016 15752 10044
rect 15252 10004 15258 10016
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 15930 10004 15936 10056
rect 15988 10004 15994 10056
rect 15841 9979 15899 9985
rect 15841 9945 15853 9979
rect 15887 9976 15899 9979
rect 16454 9979 16512 9985
rect 16454 9976 16466 9979
rect 15887 9948 16466 9976
rect 15887 9945 15899 9948
rect 15841 9939 15899 9945
rect 16454 9945 16466 9948
rect 16500 9945 16512 9979
rect 16454 9939 16512 9945
rect 1104 9818 28888 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 28888 9818
rect 1104 9744 28888 9766
rect 15746 9664 15752 9716
rect 15804 9704 15810 9716
rect 16025 9707 16083 9713
rect 16025 9704 16037 9707
rect 15804 9676 16037 9704
rect 15804 9664 15810 9676
rect 16025 9673 16037 9676
rect 16071 9673 16083 9707
rect 16025 9667 16083 9673
rect 1104 9274 28888 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 28888 9274
rect 1104 9200 28888 9222
rect 1104 8730 28888 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 28888 8730
rect 1104 8656 28888 8678
rect 28258 8576 28264 8628
rect 28316 8576 28322 8628
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8480 27951 8483
rect 28442 8480 28448 8492
rect 27939 8452 28448 8480
rect 27939 8449 27951 8452
rect 27893 8443 27951 8449
rect 28442 8440 28448 8452
rect 28500 8440 28506 8492
rect 1104 8186 28888 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 28888 8186
rect 1104 8112 28888 8134
rect 28258 8032 28264 8084
rect 28316 8072 28322 8084
rect 28353 8075 28411 8081
rect 28353 8072 28365 8075
rect 28316 8044 28365 8072
rect 28316 8032 28322 8044
rect 28353 8041 28365 8044
rect 28399 8041 28411 8075
rect 28353 8035 28411 8041
rect 1104 7642 28888 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 28888 7642
rect 1104 7568 28888 7590
rect 1104 7098 28888 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 28888 7098
rect 1104 7024 28888 7046
rect 1104 6554 28888 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 28888 6554
rect 1104 6480 28888 6502
rect 1104 6010 28888 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 28888 6010
rect 1104 5936 28888 5958
rect 1104 5466 28888 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 28888 5466
rect 1104 5392 28888 5414
rect 1104 4922 28888 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 28888 4922
rect 1104 4848 28888 4870
rect 1104 4378 28888 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 28888 3290
rect 1104 3216 28888 3238
rect 1104 2746 28888 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 28888 2746
rect 1104 2672 28888 2694
rect 5902 2592 5908 2644
rect 5960 2592 5966 2644
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 5868 2400 6101 2428
rect 5868 2388 5874 2400
rect 6089 2397 6101 2400
rect 6135 2428 6147 2431
rect 6457 2431 6515 2437
rect 6457 2428 6469 2431
rect 6135 2400 6469 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 6457 2397 6469 2400
rect 6503 2397 6515 2431
rect 6457 2391 6515 2397
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21968 2400 22017 2428
rect 21968 2388 21974 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 1104 2202 28888 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 24584 47243 24636 47252
rect 24584 47209 24593 47243
rect 24593 47209 24627 47243
rect 24627 47209 24636 47243
rect 24584 47200 24636 47209
rect 4712 47132 4764 47184
rect 22008 47064 22060 47116
rect 5448 47039 5500 47048
rect 5448 47005 5457 47039
rect 5457 47005 5491 47039
rect 5491 47005 5500 47039
rect 5448 46996 5500 47005
rect 22100 47039 22152 47048
rect 22100 47005 22109 47039
rect 22109 47005 22143 47039
rect 22143 47005 22152 47039
rect 22100 46996 22152 47005
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 10048 45500 10100 45552
rect 10876 45475 10928 45484
rect 10876 45441 10885 45475
rect 10885 45441 10919 45475
rect 10919 45441 10928 45475
rect 10876 45432 10928 45441
rect 11796 45475 11848 45484
rect 11796 45441 11805 45475
rect 11805 45441 11839 45475
rect 11839 45441 11848 45475
rect 11796 45432 11848 45441
rect 11888 45432 11940 45484
rect 11704 45364 11756 45416
rect 9956 45296 10008 45348
rect 10876 45296 10928 45348
rect 13912 45475 13964 45484
rect 13912 45441 13921 45475
rect 13921 45441 13955 45475
rect 13955 45441 13964 45475
rect 13912 45432 13964 45441
rect 14372 45364 14424 45416
rect 14740 45432 14792 45484
rect 16028 45475 16080 45484
rect 16028 45441 16037 45475
rect 16037 45441 16071 45475
rect 16071 45441 16080 45475
rect 16028 45432 16080 45441
rect 20628 45500 20680 45552
rect 19524 45432 19576 45484
rect 19984 45432 20036 45484
rect 14096 45296 14148 45348
rect 15752 45364 15804 45416
rect 18144 45364 18196 45416
rect 18420 45364 18472 45416
rect 22100 45296 22152 45348
rect 9404 45228 9456 45280
rect 11060 45228 11112 45280
rect 13820 45228 13872 45280
rect 14648 45271 14700 45280
rect 14648 45237 14657 45271
rect 14657 45237 14691 45271
rect 14691 45237 14700 45271
rect 14648 45228 14700 45237
rect 14924 45271 14976 45280
rect 14924 45237 14933 45271
rect 14933 45237 14967 45271
rect 14967 45237 14976 45271
rect 14924 45228 14976 45237
rect 16488 45228 16540 45280
rect 17500 45271 17552 45280
rect 17500 45237 17509 45271
rect 17509 45237 17543 45271
rect 17543 45237 17552 45271
rect 17500 45228 17552 45237
rect 17776 45271 17828 45280
rect 17776 45237 17785 45271
rect 17785 45237 17819 45271
rect 17819 45237 17828 45271
rect 17776 45228 17828 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 10048 45067 10100 45076
rect 10048 45033 10057 45067
rect 10057 45033 10091 45067
rect 10091 45033 10100 45067
rect 10048 45024 10100 45033
rect 7472 44863 7524 44872
rect 7472 44829 7481 44863
rect 7481 44829 7515 44863
rect 7515 44829 7524 44863
rect 7472 44820 7524 44829
rect 9496 44820 9548 44872
rect 6920 44727 6972 44736
rect 6920 44693 6929 44727
rect 6929 44693 6963 44727
rect 6963 44693 6972 44727
rect 6920 44684 6972 44693
rect 7840 44727 7892 44736
rect 7840 44693 7849 44727
rect 7849 44693 7883 44727
rect 7883 44693 7892 44727
rect 7840 44684 7892 44693
rect 9956 44752 10008 44804
rect 11704 45024 11756 45076
rect 16028 45024 16080 45076
rect 19984 45067 20036 45076
rect 19984 45033 19993 45067
rect 19993 45033 20027 45067
rect 20027 45033 20036 45067
rect 19984 45024 20036 45033
rect 11152 44888 11204 44940
rect 9220 44684 9272 44736
rect 10784 44863 10836 44872
rect 10784 44829 10793 44863
rect 10793 44829 10827 44863
rect 10827 44829 10836 44863
rect 10784 44820 10836 44829
rect 11244 44820 11296 44872
rect 11888 44820 11940 44872
rect 12532 44752 12584 44804
rect 15016 44820 15068 44872
rect 14280 44752 14332 44804
rect 14648 44752 14700 44804
rect 18420 44820 18472 44872
rect 19340 44863 19392 44872
rect 19340 44829 19349 44863
rect 19349 44829 19383 44863
rect 19383 44829 19392 44863
rect 19340 44820 19392 44829
rect 17500 44752 17552 44804
rect 12256 44684 12308 44736
rect 12440 44727 12492 44736
rect 12440 44693 12449 44727
rect 12449 44693 12483 44727
rect 12483 44693 12492 44727
rect 12440 44684 12492 44693
rect 18144 44684 18196 44736
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 10784 44480 10836 44532
rect 11244 44523 11296 44532
rect 11244 44489 11253 44523
rect 11253 44489 11287 44523
rect 11287 44489 11296 44523
rect 11244 44480 11296 44489
rect 11796 44480 11848 44532
rect 12440 44412 12492 44464
rect 4712 44387 4764 44396
rect 4712 44353 4721 44387
rect 4721 44353 4755 44387
rect 4755 44353 4764 44387
rect 4712 44344 4764 44353
rect 5632 44344 5684 44396
rect 9404 44387 9456 44396
rect 9404 44353 9413 44387
rect 9413 44353 9447 44387
rect 9447 44353 9456 44387
rect 9404 44344 9456 44353
rect 11152 44344 11204 44396
rect 4712 44140 4764 44192
rect 7196 44319 7248 44328
rect 7196 44285 7205 44319
rect 7205 44285 7239 44319
rect 7239 44285 7248 44319
rect 7196 44276 7248 44285
rect 9864 44319 9916 44328
rect 9864 44285 9873 44319
rect 9873 44285 9907 44319
rect 9907 44285 9916 44319
rect 9864 44276 9916 44285
rect 11704 44276 11756 44328
rect 11888 44319 11940 44328
rect 11888 44285 11897 44319
rect 11897 44285 11931 44319
rect 11931 44285 11940 44319
rect 11888 44276 11940 44285
rect 11520 44208 11572 44260
rect 6920 44140 6972 44192
rect 7932 44140 7984 44192
rect 8576 44183 8628 44192
rect 8576 44149 8585 44183
rect 8585 44149 8619 44183
rect 8619 44149 8628 44183
rect 8576 44140 8628 44149
rect 11796 44140 11848 44192
rect 12716 44344 12768 44396
rect 13820 44412 13872 44464
rect 13452 44387 13504 44396
rect 13452 44353 13461 44387
rect 13461 44353 13495 44387
rect 13495 44353 13504 44387
rect 13452 44344 13504 44353
rect 14096 44523 14148 44532
rect 14096 44489 14105 44523
rect 14105 44489 14139 44523
rect 14139 44489 14148 44523
rect 14096 44480 14148 44489
rect 14740 44480 14792 44532
rect 17776 44480 17828 44532
rect 16488 44412 16540 44464
rect 14280 44387 14332 44396
rect 14280 44353 14289 44387
rect 14289 44353 14323 44387
rect 14323 44353 14332 44387
rect 14280 44344 14332 44353
rect 15752 44344 15804 44396
rect 18236 44412 18288 44464
rect 18420 44412 18472 44464
rect 18052 44387 18104 44396
rect 18052 44353 18086 44387
rect 18086 44353 18104 44387
rect 14740 44208 14792 44260
rect 15568 44276 15620 44328
rect 18052 44344 18104 44353
rect 16856 44276 16908 44328
rect 20628 44387 20680 44396
rect 20628 44353 20637 44387
rect 20637 44353 20671 44387
rect 20671 44353 20680 44387
rect 20628 44344 20680 44353
rect 17684 44208 17736 44260
rect 19524 44208 19576 44260
rect 12900 44140 12952 44192
rect 14004 44140 14056 44192
rect 20076 44183 20128 44192
rect 20076 44149 20085 44183
rect 20085 44149 20119 44183
rect 20119 44149 20128 44183
rect 20076 44140 20128 44149
rect 21180 44140 21232 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 7472 43936 7524 43988
rect 11796 43936 11848 43988
rect 9864 43843 9916 43852
rect 4528 43732 4580 43784
rect 7196 43732 7248 43784
rect 9864 43809 9873 43843
rect 9873 43809 9907 43843
rect 9907 43809 9916 43843
rect 9864 43800 9916 43809
rect 12532 43868 12584 43920
rect 12900 43979 12952 43988
rect 12900 43945 12909 43979
rect 12909 43945 12943 43979
rect 12943 43945 12952 43979
rect 12900 43936 12952 43945
rect 13360 43979 13412 43988
rect 13360 43945 13369 43979
rect 13369 43945 13403 43979
rect 13403 43945 13412 43979
rect 13360 43936 13412 43945
rect 18052 43936 18104 43988
rect 20260 43979 20312 43988
rect 20260 43945 20269 43979
rect 20269 43945 20303 43979
rect 20303 43945 20312 43979
rect 20260 43936 20312 43945
rect 20628 43936 20680 43988
rect 12716 43868 12768 43920
rect 13176 43868 13228 43920
rect 14740 43868 14792 43920
rect 19340 43868 19392 43920
rect 13820 43843 13872 43852
rect 13820 43809 13829 43843
rect 13829 43809 13863 43843
rect 13863 43809 13872 43843
rect 13820 43800 13872 43809
rect 14096 43800 14148 43852
rect 14372 43800 14424 43852
rect 15016 43843 15068 43852
rect 15016 43809 15025 43843
rect 15025 43809 15059 43843
rect 15059 43809 15068 43843
rect 15016 43800 15068 43809
rect 4712 43707 4764 43716
rect 4712 43673 4746 43707
rect 4746 43673 4764 43707
rect 4712 43664 4764 43673
rect 7840 43664 7892 43716
rect 10968 43732 11020 43784
rect 11796 43775 11848 43784
rect 11796 43741 11805 43775
rect 11805 43741 11839 43775
rect 11839 43741 11848 43775
rect 11796 43732 11848 43741
rect 11888 43775 11940 43784
rect 11888 43741 11897 43775
rect 11897 43741 11931 43775
rect 11931 43741 11940 43775
rect 11888 43732 11940 43741
rect 11980 43775 12032 43784
rect 11980 43741 11989 43775
rect 11989 43741 12023 43775
rect 12023 43741 12032 43775
rect 11980 43732 12032 43741
rect 12256 43732 12308 43784
rect 9956 43664 10008 43716
rect 13544 43732 13596 43784
rect 15568 43732 15620 43784
rect 16672 43775 16724 43784
rect 16672 43741 16681 43775
rect 16681 43741 16715 43775
rect 16715 43741 16724 43775
rect 16672 43732 16724 43741
rect 16764 43775 16816 43784
rect 16764 43741 16774 43775
rect 16774 43741 16808 43775
rect 16808 43741 16816 43775
rect 16764 43732 16816 43741
rect 17132 43775 17184 43784
rect 17132 43741 17146 43775
rect 17146 43741 17180 43775
rect 17180 43741 17184 43775
rect 17132 43732 17184 43741
rect 15844 43664 15896 43716
rect 16856 43664 16908 43716
rect 16948 43707 17000 43716
rect 16948 43673 16957 43707
rect 16957 43673 16991 43707
rect 16991 43673 17000 43707
rect 16948 43664 17000 43673
rect 6460 43596 6512 43648
rect 11612 43596 11664 43648
rect 16396 43639 16448 43648
rect 16396 43605 16405 43639
rect 16405 43605 16439 43639
rect 16439 43605 16448 43639
rect 16396 43596 16448 43605
rect 16488 43596 16540 43648
rect 17224 43596 17276 43648
rect 17684 43775 17736 43784
rect 17684 43741 17693 43775
rect 17693 43741 17727 43775
rect 17727 43741 17736 43775
rect 17684 43732 17736 43741
rect 17868 43707 17920 43716
rect 17868 43673 17877 43707
rect 17877 43673 17911 43707
rect 17911 43673 17920 43707
rect 17868 43664 17920 43673
rect 19708 43775 19760 43784
rect 19708 43741 19717 43775
rect 19717 43741 19751 43775
rect 19751 43741 19760 43775
rect 19708 43732 19760 43741
rect 20628 43732 20680 43784
rect 20076 43707 20128 43716
rect 20076 43673 20085 43707
rect 20085 43673 20119 43707
rect 20119 43673 20128 43707
rect 20076 43664 20128 43673
rect 19248 43596 19300 43648
rect 21180 43639 21232 43648
rect 21180 43605 21189 43639
rect 21189 43605 21223 43639
rect 21223 43605 21232 43639
rect 21180 43596 21232 43605
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 11980 43392 12032 43444
rect 13176 43435 13228 43444
rect 13176 43401 13185 43435
rect 13185 43401 13219 43435
rect 13219 43401 13228 43435
rect 13176 43392 13228 43401
rect 15844 43435 15896 43444
rect 15844 43401 15853 43435
rect 15853 43401 15887 43435
rect 15887 43401 15896 43435
rect 15844 43392 15896 43401
rect 16764 43435 16816 43444
rect 16764 43401 16773 43435
rect 16773 43401 16807 43435
rect 16807 43401 16816 43435
rect 16764 43392 16816 43401
rect 18420 43392 18472 43444
rect 20260 43392 20312 43444
rect 11888 43324 11940 43376
rect 13912 43324 13964 43376
rect 6460 43299 6512 43308
rect 6460 43265 6469 43299
rect 6469 43265 6503 43299
rect 6503 43265 6512 43299
rect 6460 43256 6512 43265
rect 10048 43256 10100 43308
rect 11060 43256 11112 43308
rect 11612 43299 11664 43308
rect 11612 43265 11621 43299
rect 11621 43265 11655 43299
rect 11655 43265 11664 43299
rect 11612 43256 11664 43265
rect 12532 43299 12584 43308
rect 12532 43265 12541 43299
rect 12541 43265 12575 43299
rect 12575 43265 12584 43299
rect 12532 43256 12584 43265
rect 13544 43299 13596 43308
rect 13544 43265 13553 43299
rect 13553 43265 13587 43299
rect 13587 43265 13596 43299
rect 13544 43256 13596 43265
rect 14004 43299 14056 43308
rect 14004 43265 14013 43299
rect 14013 43265 14047 43299
rect 14047 43265 14056 43299
rect 14004 43256 14056 43265
rect 17040 43299 17092 43308
rect 17040 43265 17049 43299
rect 17049 43265 17083 43299
rect 17083 43265 17092 43299
rect 17040 43256 17092 43265
rect 17224 43256 17276 43308
rect 17960 43256 18012 43308
rect 18236 43299 18288 43308
rect 18236 43265 18245 43299
rect 18245 43265 18279 43299
rect 18279 43265 18288 43299
rect 18236 43256 18288 43265
rect 19340 43256 19392 43308
rect 12624 43188 12676 43240
rect 14096 43231 14148 43240
rect 14096 43197 14105 43231
rect 14105 43197 14139 43231
rect 14139 43197 14148 43231
rect 14096 43188 14148 43197
rect 15200 43231 15252 43240
rect 15200 43197 15209 43231
rect 15209 43197 15243 43231
rect 15243 43197 15252 43231
rect 15200 43188 15252 43197
rect 11980 43120 12032 43172
rect 5816 43052 5868 43104
rect 6828 43052 6880 43104
rect 11796 43052 11848 43104
rect 12440 43052 12492 43104
rect 14648 43120 14700 43172
rect 17132 43120 17184 43172
rect 17040 43052 17092 43104
rect 19708 43052 19760 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 11704 42891 11756 42900
rect 11704 42857 11713 42891
rect 11713 42857 11747 42891
rect 11747 42857 11756 42891
rect 11704 42848 11756 42857
rect 9956 42780 10008 42832
rect 16948 42848 17000 42900
rect 17960 42780 18012 42832
rect 10968 42755 11020 42764
rect 10968 42721 10977 42755
rect 10977 42721 11011 42755
rect 11011 42721 11020 42755
rect 10968 42712 11020 42721
rect 11336 42712 11388 42764
rect 12072 42755 12124 42764
rect 12072 42721 12081 42755
rect 12081 42721 12115 42755
rect 12115 42721 12124 42755
rect 12072 42712 12124 42721
rect 4712 42644 4764 42696
rect 11796 42644 11848 42696
rect 11980 42644 12032 42696
rect 12440 42687 12492 42696
rect 12440 42653 12449 42687
rect 12449 42653 12483 42687
rect 12483 42653 12492 42687
rect 12440 42644 12492 42653
rect 15200 42712 15252 42764
rect 18420 42755 18472 42764
rect 18420 42721 18429 42755
rect 18429 42721 18463 42755
rect 18463 42721 18472 42755
rect 18420 42712 18472 42721
rect 19248 42712 19300 42764
rect 19340 42755 19392 42764
rect 19340 42721 19349 42755
rect 19349 42721 19383 42755
rect 19383 42721 19392 42755
rect 19340 42712 19392 42721
rect 13544 42644 13596 42696
rect 14096 42644 14148 42696
rect 5448 42576 5500 42628
rect 11336 42619 11388 42628
rect 11336 42585 11345 42619
rect 11345 42585 11379 42619
rect 11379 42585 11388 42619
rect 11336 42576 11388 42585
rect 6460 42551 6512 42560
rect 6460 42517 6469 42551
rect 6469 42517 6503 42551
rect 6503 42517 6512 42551
rect 6460 42508 6512 42517
rect 14648 42687 14700 42696
rect 14648 42653 14657 42687
rect 14657 42653 14691 42687
rect 14691 42653 14700 42687
rect 14648 42644 14700 42653
rect 15016 42687 15068 42696
rect 15016 42653 15025 42687
rect 15025 42653 15059 42687
rect 15059 42653 15068 42687
rect 15016 42644 15068 42653
rect 15568 42576 15620 42628
rect 14740 42551 14792 42560
rect 14740 42517 14749 42551
rect 14749 42517 14783 42551
rect 14783 42517 14792 42551
rect 14740 42508 14792 42517
rect 16120 42687 16172 42696
rect 16120 42653 16129 42687
rect 16129 42653 16163 42687
rect 16163 42653 16172 42687
rect 16120 42644 16172 42653
rect 19432 42644 19484 42696
rect 16304 42619 16356 42628
rect 16304 42585 16313 42619
rect 16313 42585 16347 42619
rect 16347 42585 16356 42619
rect 16304 42576 16356 42585
rect 17040 42576 17092 42628
rect 16488 42508 16540 42560
rect 17868 42508 17920 42560
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 5448 42347 5500 42356
rect 5448 42313 5457 42347
rect 5457 42313 5491 42347
rect 5491 42313 5500 42347
rect 5448 42304 5500 42313
rect 19432 42347 19484 42356
rect 19432 42313 19441 42347
rect 19441 42313 19475 42347
rect 19475 42313 19484 42347
rect 19432 42304 19484 42313
rect 5632 42211 5684 42220
rect 5632 42177 5641 42211
rect 5641 42177 5675 42211
rect 5675 42177 5684 42211
rect 5632 42168 5684 42177
rect 5816 42211 5868 42220
rect 5816 42177 5825 42211
rect 5825 42177 5859 42211
rect 5859 42177 5868 42211
rect 5816 42168 5868 42177
rect 6460 42211 6512 42220
rect 6460 42177 6469 42211
rect 6469 42177 6503 42211
rect 6503 42177 6512 42211
rect 6460 42168 6512 42177
rect 19708 42236 19760 42288
rect 7104 42007 7156 42016
rect 7104 41973 7113 42007
rect 7113 41973 7147 42007
rect 7147 41973 7156 42007
rect 7104 41964 7156 41973
rect 20168 41964 20220 42016
rect 21180 41964 21232 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 7104 41624 7156 41676
rect 5632 41556 5684 41608
rect 12624 41556 12676 41608
rect 5540 41420 5592 41472
rect 16028 41420 16080 41472
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 6828 41216 6880 41268
rect 5448 41148 5500 41200
rect 6644 41148 6696 41200
rect 4712 41123 4764 41132
rect 4712 41089 4721 41123
rect 4721 41089 4755 41123
rect 4755 41089 4764 41123
rect 4712 41080 4764 41089
rect 5540 41080 5592 41132
rect 7196 41148 7248 41200
rect 7932 41080 7984 41132
rect 7472 40876 7524 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 6828 40715 6880 40724
rect 6828 40681 6837 40715
rect 6837 40681 6871 40715
rect 6871 40681 6880 40715
rect 6828 40672 6880 40681
rect 7748 40672 7800 40724
rect 8576 40672 8628 40724
rect 9496 40715 9548 40724
rect 9496 40681 9505 40715
rect 9505 40681 9539 40715
rect 9539 40681 9548 40715
rect 9496 40672 9548 40681
rect 10692 40672 10744 40724
rect 16304 40672 16356 40724
rect 10876 40604 10928 40656
rect 7656 40536 7708 40588
rect 7840 40536 7892 40588
rect 7932 40579 7984 40588
rect 7932 40545 7941 40579
rect 7941 40545 7975 40579
rect 7975 40545 7984 40579
rect 7932 40536 7984 40545
rect 5632 40468 5684 40520
rect 6644 40511 6696 40520
rect 6644 40477 6653 40511
rect 6653 40477 6687 40511
rect 6687 40477 6696 40511
rect 6644 40468 6696 40477
rect 7104 40468 7156 40520
rect 10968 40468 11020 40520
rect 16028 40511 16080 40520
rect 16028 40477 16037 40511
rect 16037 40477 16071 40511
rect 16071 40477 16080 40511
rect 16028 40468 16080 40477
rect 7288 40400 7340 40452
rect 5908 40375 5960 40384
rect 5908 40341 5917 40375
rect 5917 40341 5951 40375
rect 5951 40341 5960 40375
rect 5908 40332 5960 40341
rect 15844 40443 15896 40452
rect 15844 40409 15853 40443
rect 15853 40409 15887 40443
rect 15887 40409 15896 40443
rect 15844 40400 15896 40409
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 7656 40171 7708 40180
rect 7656 40137 7665 40171
rect 7665 40137 7699 40171
rect 7699 40137 7708 40171
rect 7656 40128 7708 40137
rect 7840 40128 7892 40180
rect 10968 40171 11020 40180
rect 10968 40137 10977 40171
rect 10977 40137 11011 40171
rect 11011 40137 11020 40171
rect 10968 40128 11020 40137
rect 11612 40171 11664 40180
rect 11612 40137 11621 40171
rect 11621 40137 11655 40171
rect 11655 40137 11664 40171
rect 11612 40128 11664 40137
rect 16212 40128 16264 40180
rect 16672 40128 16724 40180
rect 8024 39992 8076 40044
rect 8208 40035 8260 40044
rect 8208 40001 8242 40035
rect 8242 40001 8260 40035
rect 8208 39992 8260 40001
rect 9680 39992 9732 40044
rect 11244 39992 11296 40044
rect 7012 39967 7064 39976
rect 7012 39933 7021 39967
rect 7021 39933 7055 39967
rect 7055 39933 7064 39967
rect 7012 39924 7064 39933
rect 11428 39924 11480 39976
rect 11152 39856 11204 39908
rect 13176 39924 13228 39976
rect 15292 39992 15344 40044
rect 15568 40035 15620 40044
rect 15568 40001 15577 40035
rect 15577 40001 15611 40035
rect 15611 40001 15620 40035
rect 15568 39992 15620 40001
rect 15200 39924 15252 39976
rect 17868 39924 17920 39976
rect 15752 39856 15804 39908
rect 15660 39788 15712 39840
rect 16396 39831 16448 39840
rect 16396 39797 16405 39831
rect 16405 39797 16439 39831
rect 16439 39797 16448 39831
rect 16396 39788 16448 39797
rect 18420 39788 18472 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 7012 39627 7064 39636
rect 7012 39593 7021 39627
rect 7021 39593 7055 39627
rect 7055 39593 7064 39627
rect 7012 39584 7064 39593
rect 8208 39584 8260 39636
rect 9680 39584 9732 39636
rect 16120 39584 16172 39636
rect 5540 39448 5592 39500
rect 7656 39448 7708 39500
rect 15292 39516 15344 39568
rect 10876 39448 10928 39500
rect 5908 39423 5960 39432
rect 5908 39389 5942 39423
rect 5942 39389 5960 39423
rect 5908 39380 5960 39389
rect 9220 39423 9272 39432
rect 9220 39389 9229 39423
rect 9229 39389 9263 39423
rect 9263 39389 9272 39423
rect 9220 39380 9272 39389
rect 7288 39312 7340 39364
rect 7840 39312 7892 39364
rect 10784 39423 10836 39432
rect 10784 39389 10793 39423
rect 10793 39389 10827 39423
rect 10827 39389 10836 39423
rect 10784 39380 10836 39389
rect 11428 39448 11480 39500
rect 12072 39491 12124 39500
rect 12072 39457 12081 39491
rect 12081 39457 12115 39491
rect 12115 39457 12124 39491
rect 12072 39448 12124 39457
rect 10692 39312 10744 39364
rect 8668 39287 8720 39296
rect 8668 39253 8677 39287
rect 8677 39253 8711 39287
rect 8711 39253 8720 39287
rect 8668 39244 8720 39253
rect 9036 39244 9088 39296
rect 13636 39380 13688 39432
rect 19524 39448 19576 39500
rect 15476 39423 15528 39432
rect 15476 39389 15486 39423
rect 15486 39389 15520 39423
rect 15520 39389 15528 39423
rect 15476 39380 15528 39389
rect 15660 39423 15712 39432
rect 15660 39389 15669 39423
rect 15669 39389 15703 39423
rect 15703 39389 15712 39423
rect 15660 39380 15712 39389
rect 15844 39423 15896 39432
rect 15844 39389 15858 39423
rect 15858 39389 15892 39423
rect 15892 39389 15896 39423
rect 15844 39380 15896 39389
rect 15200 39312 15252 39364
rect 15568 39312 15620 39364
rect 16028 39312 16080 39364
rect 16396 39423 16448 39432
rect 16396 39389 16405 39423
rect 16405 39389 16439 39423
rect 16439 39389 16448 39423
rect 16396 39380 16448 39389
rect 18420 39423 18472 39432
rect 18420 39389 18429 39423
rect 18429 39389 18463 39423
rect 18463 39389 18472 39423
rect 18420 39380 18472 39389
rect 18696 39423 18748 39432
rect 18696 39389 18705 39423
rect 18705 39389 18739 39423
rect 18739 39389 18748 39423
rect 18696 39380 18748 39389
rect 16488 39312 16540 39364
rect 16856 39244 16908 39296
rect 19156 39244 19208 39296
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 7748 39083 7800 39092
rect 7748 39049 7757 39083
rect 7757 39049 7791 39083
rect 7791 39049 7800 39083
rect 7748 39040 7800 39049
rect 10784 39040 10836 39092
rect 13176 39083 13228 39092
rect 13176 39049 13185 39083
rect 13185 39049 13219 39083
rect 13219 39049 13228 39083
rect 13176 39040 13228 39049
rect 17868 39083 17920 39092
rect 17868 39049 17877 39083
rect 17877 39049 17911 39083
rect 17911 39049 17920 39083
rect 17868 39040 17920 39049
rect 18696 39040 18748 39092
rect 8208 38972 8260 39024
rect 8668 39015 8720 39024
rect 8668 38981 8702 39015
rect 8702 38981 8720 39015
rect 8668 38972 8720 38981
rect 7472 38947 7524 38956
rect 7472 38913 7481 38947
rect 7481 38913 7515 38947
rect 7515 38913 7524 38947
rect 7472 38904 7524 38913
rect 7840 38947 7892 38956
rect 7840 38913 7849 38947
rect 7849 38913 7883 38947
rect 7883 38913 7892 38947
rect 7840 38904 7892 38913
rect 8024 38904 8076 38956
rect 9036 38904 9088 38956
rect 10508 38904 10560 38956
rect 11060 38904 11112 38956
rect 12072 38904 12124 38956
rect 12716 38904 12768 38956
rect 13636 38947 13688 38956
rect 13636 38913 13645 38947
rect 13645 38913 13679 38947
rect 13679 38913 13688 38947
rect 13636 38904 13688 38913
rect 13912 38947 13964 38956
rect 13912 38913 13921 38947
rect 13921 38913 13955 38947
rect 13955 38913 13964 38947
rect 13912 38904 13964 38913
rect 14096 38947 14148 38956
rect 14096 38913 14105 38947
rect 14105 38913 14139 38947
rect 14139 38913 14148 38947
rect 14096 38904 14148 38913
rect 15844 38947 15896 38956
rect 15844 38913 15853 38947
rect 15853 38913 15887 38947
rect 15887 38913 15896 38947
rect 15844 38904 15896 38913
rect 10600 38879 10652 38888
rect 10600 38845 10609 38879
rect 10609 38845 10643 38879
rect 10643 38845 10652 38879
rect 10600 38836 10652 38845
rect 11888 38836 11940 38888
rect 12808 38879 12860 38888
rect 12808 38845 12817 38879
rect 12817 38845 12851 38879
rect 12851 38845 12860 38879
rect 12808 38836 12860 38845
rect 13176 38836 13228 38888
rect 15568 38836 15620 38888
rect 16304 38904 16356 38956
rect 16856 38947 16908 38956
rect 16856 38913 16865 38947
rect 16865 38913 16899 38947
rect 16899 38913 16908 38947
rect 16856 38904 16908 38913
rect 19156 38904 19208 38956
rect 19524 38947 19576 38956
rect 19524 38913 19533 38947
rect 19533 38913 19567 38947
rect 19567 38913 19576 38947
rect 19524 38904 19576 38913
rect 19800 38972 19852 39024
rect 19984 38947 20036 38956
rect 19984 38913 19993 38947
rect 19993 38913 20027 38947
rect 20027 38913 20036 38947
rect 19984 38904 20036 38913
rect 20168 38947 20220 38956
rect 20168 38913 20177 38947
rect 20177 38913 20211 38947
rect 20211 38913 20220 38947
rect 20168 38904 20220 38913
rect 18144 38836 18196 38888
rect 12532 38768 12584 38820
rect 10048 38743 10100 38752
rect 10048 38709 10057 38743
rect 10057 38709 10091 38743
rect 10091 38709 10100 38743
rect 10048 38700 10100 38709
rect 11796 38700 11848 38752
rect 12164 38700 12216 38752
rect 12348 38700 12400 38752
rect 14004 38743 14056 38752
rect 14004 38709 14013 38743
rect 14013 38709 14047 38743
rect 14047 38709 14056 38743
rect 14004 38700 14056 38709
rect 15384 38700 15436 38752
rect 17592 38700 17644 38752
rect 18236 38700 18288 38752
rect 19524 38743 19576 38752
rect 19524 38709 19533 38743
rect 19533 38709 19567 38743
rect 19567 38709 19576 38743
rect 19524 38700 19576 38709
rect 23112 38700 23164 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 9036 38539 9088 38548
rect 9036 38505 9045 38539
rect 9045 38505 9079 38539
rect 9079 38505 9088 38539
rect 9036 38496 9088 38505
rect 9220 38496 9272 38548
rect 9588 38496 9640 38548
rect 11060 38471 11112 38480
rect 11060 38437 11069 38471
rect 11069 38437 11103 38471
rect 11103 38437 11112 38471
rect 11060 38428 11112 38437
rect 10048 38360 10100 38412
rect 1216 38292 1268 38344
rect 7288 38292 7340 38344
rect 1676 38199 1728 38208
rect 1676 38165 1685 38199
rect 1685 38165 1719 38199
rect 1719 38165 1728 38199
rect 1676 38156 1728 38165
rect 10324 38199 10376 38208
rect 10324 38165 10333 38199
rect 10333 38165 10367 38199
rect 10367 38165 10376 38199
rect 10324 38156 10376 38165
rect 10508 38335 10560 38344
rect 10508 38301 10517 38335
rect 10517 38301 10551 38335
rect 10551 38301 10560 38335
rect 10508 38292 10560 38301
rect 12716 38496 12768 38548
rect 16856 38496 16908 38548
rect 15568 38471 15620 38480
rect 15568 38437 15577 38471
rect 15577 38437 15611 38471
rect 15611 38437 15620 38471
rect 15568 38428 15620 38437
rect 19340 38496 19392 38548
rect 19984 38496 20036 38548
rect 15292 38360 15344 38412
rect 16488 38360 16540 38412
rect 16856 38360 16908 38412
rect 17592 38403 17644 38412
rect 17592 38369 17601 38403
rect 17601 38369 17635 38403
rect 17635 38369 17644 38403
rect 17592 38360 17644 38369
rect 12164 38335 12216 38344
rect 12164 38301 12182 38335
rect 12182 38301 12216 38335
rect 12164 38292 12216 38301
rect 12348 38224 12400 38276
rect 12256 38156 12308 38208
rect 12900 38292 12952 38344
rect 13084 38335 13136 38344
rect 13084 38301 13093 38335
rect 13093 38301 13127 38335
rect 13127 38301 13136 38335
rect 13084 38292 13136 38301
rect 13176 38335 13228 38344
rect 13176 38301 13185 38335
rect 13185 38301 13219 38335
rect 13219 38301 13228 38335
rect 13176 38292 13228 38301
rect 14004 38292 14056 38344
rect 15844 38335 15896 38344
rect 15844 38301 15853 38335
rect 15853 38301 15887 38335
rect 15887 38301 15896 38335
rect 15844 38292 15896 38301
rect 16212 38292 16264 38344
rect 16120 38224 16172 38276
rect 16764 38292 16816 38344
rect 19800 38292 19852 38344
rect 16580 38224 16632 38276
rect 18604 38224 18656 38276
rect 15660 38156 15712 38208
rect 17776 38156 17828 38208
rect 19892 38156 19944 38208
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 9036 37952 9088 38004
rect 10508 37952 10560 38004
rect 12808 37952 12860 38004
rect 13084 37952 13136 38004
rect 14096 37952 14148 38004
rect 1676 37816 1728 37868
rect 5448 37884 5500 37936
rect 5356 37748 5408 37800
rect 9588 37884 9640 37936
rect 9036 37816 9088 37868
rect 11152 37816 11204 37868
rect 11244 37859 11296 37868
rect 11244 37825 11253 37859
rect 11253 37825 11287 37859
rect 11287 37825 11296 37859
rect 11244 37816 11296 37825
rect 12992 37884 13044 37936
rect 14740 37884 14792 37936
rect 15384 37927 15436 37936
rect 15384 37893 15393 37927
rect 15393 37893 15427 37927
rect 15427 37893 15436 37927
rect 15384 37884 15436 37893
rect 16120 37927 16172 37936
rect 16120 37893 16129 37927
rect 16129 37893 16163 37927
rect 16163 37893 16172 37927
rect 16120 37884 16172 37893
rect 11796 37859 11848 37868
rect 11796 37825 11805 37859
rect 11805 37825 11839 37859
rect 11839 37825 11848 37859
rect 11796 37816 11848 37825
rect 11888 37859 11940 37868
rect 11888 37825 11897 37859
rect 11897 37825 11931 37859
rect 11931 37825 11940 37859
rect 11888 37816 11940 37825
rect 12348 37816 12400 37868
rect 14188 37859 14240 37868
rect 14188 37825 14197 37859
rect 14197 37825 14231 37859
rect 14231 37825 14240 37859
rect 14188 37816 14240 37825
rect 14464 37859 14516 37868
rect 14464 37825 14473 37859
rect 14473 37825 14507 37859
rect 14507 37825 14516 37859
rect 14464 37816 14516 37825
rect 15200 37859 15252 37868
rect 15200 37825 15204 37859
rect 15204 37825 15238 37859
rect 15238 37825 15252 37859
rect 7012 37748 7064 37800
rect 4804 37612 4856 37664
rect 7288 37680 7340 37732
rect 8024 37748 8076 37800
rect 12624 37748 12676 37800
rect 15200 37816 15252 37825
rect 15568 37859 15620 37868
rect 15568 37825 15576 37859
rect 15576 37825 15610 37859
rect 15610 37825 15620 37859
rect 15568 37816 15620 37825
rect 15660 37859 15712 37868
rect 15660 37825 15669 37859
rect 15669 37825 15703 37859
rect 15703 37825 15712 37859
rect 15660 37816 15712 37825
rect 18604 37995 18656 38004
rect 18604 37961 18613 37995
rect 18613 37961 18647 37995
rect 18647 37961 18656 37995
rect 18604 37952 18656 37961
rect 19432 37952 19484 38004
rect 15936 37748 15988 37800
rect 17316 37791 17368 37800
rect 17316 37757 17325 37791
rect 17325 37757 17359 37791
rect 17359 37757 17368 37791
rect 17316 37748 17368 37757
rect 17868 37748 17920 37800
rect 18420 37748 18472 37800
rect 19892 37791 19944 37800
rect 19892 37757 19901 37791
rect 19901 37757 19935 37791
rect 19935 37757 19944 37791
rect 19892 37748 19944 37757
rect 15476 37680 15528 37732
rect 5632 37655 5684 37664
rect 5632 37621 5641 37655
rect 5641 37621 5675 37655
rect 5675 37621 5684 37655
rect 5632 37612 5684 37621
rect 10508 37612 10560 37664
rect 17684 37655 17736 37664
rect 17684 37621 17693 37655
rect 17693 37621 17727 37655
rect 17727 37621 17736 37655
rect 17684 37612 17736 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 11152 37408 11204 37460
rect 12440 37408 12492 37460
rect 12900 37408 12952 37460
rect 14188 37408 14240 37460
rect 16488 37408 16540 37460
rect 9036 37315 9088 37324
rect 9036 37281 9045 37315
rect 9045 37281 9079 37315
rect 9079 37281 9088 37315
rect 9036 37272 9088 37281
rect 11428 37340 11480 37392
rect 11060 37272 11112 37324
rect 7012 37247 7064 37256
rect 7012 37213 7021 37247
rect 7021 37213 7055 37247
rect 7055 37213 7064 37247
rect 7012 37204 7064 37213
rect 10324 37204 10376 37256
rect 5264 37179 5316 37188
rect 5264 37145 5298 37179
rect 5298 37145 5316 37179
rect 5264 37136 5316 37145
rect 5448 37136 5500 37188
rect 6368 37111 6420 37120
rect 6368 37077 6377 37111
rect 6377 37077 6411 37111
rect 6411 37077 6420 37111
rect 6368 37068 6420 37077
rect 13912 37340 13964 37392
rect 12348 37272 12400 37324
rect 12808 37315 12860 37324
rect 12808 37281 12817 37315
rect 12817 37281 12851 37315
rect 12851 37281 12860 37315
rect 12808 37272 12860 37281
rect 12900 37247 12952 37256
rect 12900 37213 12909 37247
rect 12909 37213 12943 37247
rect 12943 37213 12952 37247
rect 12900 37204 12952 37213
rect 13544 37247 13596 37256
rect 13544 37213 13553 37247
rect 13553 37213 13587 37247
rect 13587 37213 13596 37247
rect 13544 37204 13596 37213
rect 14648 37247 14700 37256
rect 14648 37213 14657 37247
rect 14657 37213 14691 37247
rect 14691 37213 14700 37247
rect 14648 37204 14700 37213
rect 14740 37247 14792 37256
rect 14740 37213 14749 37247
rect 14749 37213 14783 37247
rect 14783 37213 14792 37247
rect 14740 37204 14792 37213
rect 17592 37315 17644 37324
rect 17592 37281 17601 37315
rect 17601 37281 17635 37315
rect 17635 37281 17644 37315
rect 17592 37272 17644 37281
rect 17868 37408 17920 37460
rect 18420 37451 18472 37460
rect 18420 37417 18429 37451
rect 18429 37417 18463 37451
rect 18463 37417 18472 37451
rect 18420 37408 18472 37417
rect 19892 37272 19944 37324
rect 14464 37136 14516 37188
rect 17684 37204 17736 37256
rect 19524 37204 19576 37256
rect 15936 37179 15988 37188
rect 15936 37145 15945 37179
rect 15945 37145 15979 37179
rect 15979 37145 15988 37179
rect 15936 37136 15988 37145
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 5264 36864 5316 36916
rect 12900 36907 12952 36916
rect 12900 36873 12909 36907
rect 12909 36873 12943 36907
rect 12943 36873 12952 36907
rect 12900 36864 12952 36873
rect 14648 36864 14700 36916
rect 15200 36864 15252 36916
rect 12348 36796 12400 36848
rect 4804 36728 4856 36780
rect 5632 36728 5684 36780
rect 11244 36728 11296 36780
rect 11704 36728 11756 36780
rect 12440 36771 12492 36780
rect 12440 36737 12449 36771
rect 12449 36737 12483 36771
rect 12483 36737 12492 36771
rect 12440 36728 12492 36737
rect 16580 36864 16632 36916
rect 17868 36864 17920 36916
rect 16212 36796 16264 36848
rect 15936 36771 15988 36780
rect 15936 36737 15945 36771
rect 15945 36737 15979 36771
rect 15979 36737 15988 36771
rect 15936 36728 15988 36737
rect 6368 36660 6420 36712
rect 12532 36592 12584 36644
rect 17316 36592 17368 36644
rect 5632 36524 5684 36576
rect 16028 36524 16080 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 5356 36116 5408 36168
rect 6460 36116 6512 36168
rect 5540 36091 5592 36100
rect 5540 36057 5574 36091
rect 5574 36057 5592 36091
rect 5540 36048 5592 36057
rect 4804 35980 4856 36032
rect 6092 35980 6144 36032
rect 6920 36023 6972 36032
rect 6920 35989 6929 36023
rect 6929 35989 6963 36023
rect 6963 35989 6972 36023
rect 6920 35980 6972 35989
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 5540 35776 5592 35828
rect 6460 35819 6512 35828
rect 6460 35785 6469 35819
rect 6469 35785 6503 35819
rect 6503 35785 6512 35819
rect 6460 35776 6512 35785
rect 16212 35819 16264 35828
rect 16212 35785 16221 35819
rect 16221 35785 16255 35819
rect 16255 35785 16264 35819
rect 16212 35776 16264 35785
rect 16764 35819 16816 35828
rect 16764 35785 16773 35819
rect 16773 35785 16807 35819
rect 16807 35785 16816 35819
rect 16764 35776 16816 35785
rect 4804 35640 4856 35692
rect 5632 35708 5684 35760
rect 4988 35683 5040 35692
rect 4988 35649 4997 35683
rect 4997 35649 5031 35683
rect 5031 35649 5040 35683
rect 4988 35640 5040 35649
rect 5540 35640 5592 35692
rect 6920 35708 6972 35760
rect 6092 35615 6144 35624
rect 6092 35581 6101 35615
rect 6101 35581 6135 35615
rect 6135 35581 6144 35615
rect 6092 35572 6144 35581
rect 6552 35572 6604 35624
rect 8024 35640 8076 35692
rect 16304 35683 16356 35692
rect 16304 35649 16313 35683
rect 16313 35649 16347 35683
rect 16347 35649 16356 35683
rect 16304 35640 16356 35649
rect 5264 35436 5316 35488
rect 5540 35436 5592 35488
rect 6092 35436 6144 35488
rect 6920 35436 6972 35488
rect 15108 35436 15160 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 5356 35275 5408 35284
rect 5356 35241 5365 35275
rect 5365 35241 5399 35275
rect 5399 35241 5408 35275
rect 5356 35232 5408 35241
rect 6368 35164 6420 35216
rect 5540 35096 5592 35148
rect 5448 34892 5500 34944
rect 5816 35003 5868 35012
rect 5816 34969 5825 35003
rect 5825 34969 5859 35003
rect 5859 34969 5868 35003
rect 5816 34960 5868 34969
rect 5908 35003 5960 35012
rect 5908 34969 5917 35003
rect 5917 34969 5951 35003
rect 5951 34969 5960 35003
rect 5908 34960 5960 34969
rect 11704 35275 11756 35284
rect 11704 35241 11713 35275
rect 11713 35241 11747 35275
rect 11747 35241 11756 35275
rect 11704 35232 11756 35241
rect 16396 35232 16448 35284
rect 6828 35164 6880 35216
rect 16764 35164 16816 35216
rect 17592 35164 17644 35216
rect 7012 35028 7064 35080
rect 12992 35096 13044 35148
rect 9404 35071 9456 35080
rect 9404 35037 9413 35071
rect 9413 35037 9447 35071
rect 9447 35037 9456 35071
rect 9404 35028 9456 35037
rect 11888 35071 11940 35080
rect 11888 35037 11897 35071
rect 11897 35037 11931 35071
rect 11931 35037 11940 35071
rect 11888 35028 11940 35037
rect 12072 35028 12124 35080
rect 16580 35071 16632 35080
rect 16580 35037 16589 35071
rect 16589 35037 16623 35071
rect 16623 35037 16632 35071
rect 16580 35028 16632 35037
rect 9128 34960 9180 35012
rect 6184 34935 6236 34944
rect 6184 34901 6193 34935
rect 6193 34901 6227 34935
rect 6227 34901 6236 34935
rect 6184 34892 6236 34901
rect 6460 34892 6512 34944
rect 6552 34892 6604 34944
rect 6920 34892 6972 34944
rect 12348 34892 12400 34944
rect 14924 34892 14976 34944
rect 16304 34892 16356 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 5724 34688 5776 34740
rect 6828 34688 6880 34740
rect 7012 34731 7064 34740
rect 7012 34697 7021 34731
rect 7021 34697 7055 34731
rect 7055 34697 7064 34731
rect 7012 34688 7064 34697
rect 6184 34620 6236 34672
rect 5264 34595 5316 34604
rect 5264 34561 5273 34595
rect 5273 34561 5307 34595
rect 5307 34561 5316 34595
rect 5264 34552 5316 34561
rect 5632 34552 5684 34604
rect 6736 34595 6788 34604
rect 6736 34561 6745 34595
rect 6745 34561 6779 34595
rect 6779 34561 6788 34595
rect 6736 34552 6788 34561
rect 6828 34595 6880 34604
rect 6828 34561 6837 34595
rect 6837 34561 6871 34595
rect 6871 34561 6880 34595
rect 6828 34552 6880 34561
rect 10600 34688 10652 34740
rect 12992 34731 13044 34740
rect 12992 34697 13001 34731
rect 13001 34697 13035 34731
rect 13035 34697 13044 34731
rect 12992 34688 13044 34697
rect 14740 34688 14792 34740
rect 16212 34731 16264 34740
rect 10508 34663 10560 34672
rect 10508 34629 10517 34663
rect 10517 34629 10551 34663
rect 10551 34629 10560 34663
rect 10508 34620 10560 34629
rect 9864 34595 9916 34604
rect 9864 34561 9873 34595
rect 9873 34561 9907 34595
rect 9907 34561 9916 34595
rect 9864 34552 9916 34561
rect 10140 34552 10192 34604
rect 5724 34484 5776 34536
rect 6460 34527 6512 34536
rect 6460 34493 6469 34527
rect 6469 34493 6503 34527
rect 6503 34493 6512 34527
rect 6460 34484 6512 34493
rect 9404 34527 9456 34536
rect 9404 34493 9413 34527
rect 9413 34493 9447 34527
rect 9447 34493 9456 34527
rect 9404 34484 9456 34493
rect 9680 34484 9732 34536
rect 9956 34527 10008 34536
rect 9956 34493 9965 34527
rect 9965 34493 9999 34527
rect 9999 34493 10008 34527
rect 9956 34484 10008 34493
rect 10876 34620 10928 34672
rect 12808 34620 12860 34672
rect 16212 34697 16221 34731
rect 16221 34697 16255 34731
rect 16255 34697 16264 34731
rect 16212 34688 16264 34697
rect 10784 34552 10836 34604
rect 12256 34595 12308 34604
rect 12256 34561 12265 34595
rect 12265 34561 12299 34595
rect 12299 34561 12308 34595
rect 12256 34552 12308 34561
rect 14188 34595 14240 34604
rect 14188 34561 14197 34595
rect 14197 34561 14231 34595
rect 14231 34561 14240 34595
rect 14188 34552 14240 34561
rect 14648 34552 14700 34604
rect 15384 34620 15436 34672
rect 16396 34620 16448 34672
rect 14924 34595 14976 34604
rect 14924 34561 14933 34595
rect 14933 34561 14967 34595
rect 14967 34561 14976 34595
rect 14924 34552 14976 34561
rect 15108 34595 15160 34604
rect 15108 34561 15117 34595
rect 15117 34561 15151 34595
rect 15151 34561 15160 34595
rect 15108 34552 15160 34561
rect 15568 34595 15620 34604
rect 15568 34561 15577 34595
rect 15577 34561 15611 34595
rect 15611 34561 15620 34595
rect 15568 34552 15620 34561
rect 11244 34484 11296 34536
rect 19432 34527 19484 34536
rect 19432 34493 19441 34527
rect 19441 34493 19475 34527
rect 19475 34493 19484 34527
rect 19432 34484 19484 34493
rect 9036 34416 9088 34468
rect 15384 34416 15436 34468
rect 4896 34391 4948 34400
rect 4896 34357 4905 34391
rect 4905 34357 4939 34391
rect 4939 34357 4948 34391
rect 4896 34348 4948 34357
rect 7932 34391 7984 34400
rect 7932 34357 7941 34391
rect 7941 34357 7975 34391
rect 7975 34357 7984 34391
rect 7932 34348 7984 34357
rect 15292 34391 15344 34400
rect 15292 34357 15301 34391
rect 15301 34357 15335 34391
rect 15335 34357 15344 34391
rect 15292 34348 15344 34357
rect 17868 34348 17920 34400
rect 18788 34391 18840 34400
rect 18788 34357 18797 34391
rect 18797 34357 18831 34391
rect 18831 34357 18840 34391
rect 18788 34348 18840 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 5632 34187 5684 34196
rect 5632 34153 5641 34187
rect 5641 34153 5675 34187
rect 5675 34153 5684 34187
rect 5632 34144 5684 34153
rect 5816 34144 5868 34196
rect 9680 34144 9732 34196
rect 9956 34144 10008 34196
rect 12348 34144 12400 34196
rect 12624 34076 12676 34128
rect 6920 33983 6972 33992
rect 6920 33949 6929 33983
rect 6929 33949 6963 33983
rect 6963 33949 6972 33983
rect 6920 33940 6972 33949
rect 7196 33940 7248 33992
rect 9128 33940 9180 33992
rect 10692 33983 10744 33992
rect 10692 33949 10701 33983
rect 10701 33949 10735 33983
rect 10735 33949 10744 33983
rect 10692 33940 10744 33949
rect 11244 33983 11296 33992
rect 11244 33949 11253 33983
rect 11253 33949 11287 33983
rect 11287 33949 11296 33983
rect 11244 33940 11296 33949
rect 11520 33983 11572 33992
rect 11520 33949 11529 33983
rect 11529 33949 11563 33983
rect 11563 33949 11572 33983
rect 11520 33940 11572 33949
rect 12532 33983 12584 33992
rect 12532 33949 12541 33983
rect 12541 33949 12575 33983
rect 12575 33949 12584 33983
rect 12532 33940 12584 33949
rect 15844 34144 15896 34196
rect 16580 34144 16632 34196
rect 18788 34144 18840 34196
rect 17592 34008 17644 34060
rect 4896 33872 4948 33924
rect 7932 33872 7984 33924
rect 12716 33983 12768 33992
rect 12716 33949 12725 33983
rect 12725 33949 12759 33983
rect 12759 33949 12768 33983
rect 12716 33940 12768 33949
rect 12992 33940 13044 33992
rect 14372 33940 14424 33992
rect 14648 33983 14700 33992
rect 14648 33949 14657 33983
rect 14657 33949 14691 33983
rect 14691 33949 14700 33983
rect 14648 33940 14700 33949
rect 15016 33940 15068 33992
rect 17684 33940 17736 33992
rect 19156 33940 19208 33992
rect 22192 33983 22244 33992
rect 22192 33949 22201 33983
rect 22201 33949 22235 33983
rect 22235 33949 22244 33983
rect 22192 33940 22244 33949
rect 25044 33983 25096 33992
rect 25044 33949 25053 33983
rect 25053 33949 25087 33983
rect 25087 33949 25096 33983
rect 25044 33940 25096 33949
rect 12808 33872 12860 33924
rect 15292 33872 15344 33924
rect 17500 33915 17552 33924
rect 17500 33881 17509 33915
rect 17509 33881 17543 33915
rect 17543 33881 17552 33915
rect 17500 33872 17552 33881
rect 12440 33804 12492 33856
rect 13820 33847 13872 33856
rect 13820 33813 13829 33847
rect 13829 33813 13863 33847
rect 13863 33813 13872 33847
rect 13820 33804 13872 33813
rect 14556 33847 14608 33856
rect 14556 33813 14565 33847
rect 14565 33813 14599 33847
rect 14599 33813 14608 33847
rect 14556 33804 14608 33813
rect 18052 33804 18104 33856
rect 19340 33804 19392 33856
rect 19984 33847 20036 33856
rect 19984 33813 19993 33847
rect 19993 33813 20027 33847
rect 20027 33813 20036 33847
rect 19984 33804 20036 33813
rect 21548 33804 21600 33856
rect 24492 33847 24544 33856
rect 24492 33813 24501 33847
rect 24501 33813 24535 33847
rect 24535 33813 24544 33847
rect 24492 33804 24544 33813
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 9036 33600 9088 33652
rect 9956 33600 10008 33652
rect 11520 33600 11572 33652
rect 15568 33600 15620 33652
rect 19156 33643 19208 33652
rect 19156 33609 19165 33643
rect 19165 33609 19199 33643
rect 19199 33609 19208 33643
rect 19156 33600 19208 33609
rect 19432 33600 19484 33652
rect 10140 33575 10192 33584
rect 10140 33541 10174 33575
rect 10174 33541 10192 33575
rect 10140 33532 10192 33541
rect 11704 33575 11756 33584
rect 11704 33541 11713 33575
rect 11713 33541 11747 33575
rect 11747 33541 11756 33575
rect 11704 33532 11756 33541
rect 11888 33532 11940 33584
rect 14556 33532 14608 33584
rect 5632 33464 5684 33516
rect 9680 33507 9732 33516
rect 9680 33473 9689 33507
rect 9689 33473 9723 33507
rect 9723 33473 9732 33507
rect 9680 33464 9732 33473
rect 9864 33464 9916 33516
rect 12440 33507 12492 33516
rect 12440 33473 12449 33507
rect 12449 33473 12483 33507
rect 12483 33473 12492 33507
rect 12440 33464 12492 33473
rect 14188 33464 14240 33516
rect 14464 33507 14516 33516
rect 14464 33473 14473 33507
rect 14473 33473 14507 33507
rect 14507 33473 14516 33507
rect 14464 33464 14516 33473
rect 15016 33507 15068 33516
rect 15016 33473 15025 33507
rect 15025 33473 15059 33507
rect 15059 33473 15068 33507
rect 15016 33464 15068 33473
rect 17592 33464 17644 33516
rect 17868 33532 17920 33584
rect 18052 33507 18104 33516
rect 18052 33473 18086 33507
rect 18086 33473 18104 33507
rect 18052 33464 18104 33473
rect 10600 33439 10652 33448
rect 10600 33405 10609 33439
rect 10609 33405 10643 33439
rect 10643 33405 10652 33439
rect 10600 33396 10652 33405
rect 13820 33396 13872 33448
rect 14280 33396 14332 33448
rect 19984 33464 20036 33516
rect 19708 33396 19760 33448
rect 12072 33371 12124 33380
rect 12072 33337 12081 33371
rect 12081 33337 12115 33371
rect 12115 33337 12124 33371
rect 12072 33328 12124 33337
rect 12532 33328 12584 33380
rect 14096 33328 14148 33380
rect 5540 33260 5592 33312
rect 7196 33260 7248 33312
rect 11060 33260 11112 33312
rect 11888 33260 11940 33312
rect 13084 33303 13136 33312
rect 13084 33269 13093 33303
rect 13093 33269 13127 33303
rect 13127 33269 13136 33303
rect 13084 33260 13136 33269
rect 13912 33260 13964 33312
rect 21548 33507 21600 33516
rect 21548 33473 21557 33507
rect 21557 33473 21591 33507
rect 21591 33473 21600 33507
rect 21548 33464 21600 33473
rect 23756 33507 23808 33516
rect 23756 33473 23765 33507
rect 23765 33473 23799 33507
rect 23799 33473 23808 33507
rect 23756 33464 23808 33473
rect 24492 33532 24544 33584
rect 23572 33328 23624 33380
rect 23296 33303 23348 33312
rect 23296 33269 23305 33303
rect 23305 33269 23339 33303
rect 23339 33269 23348 33303
rect 23296 33260 23348 33269
rect 23664 33303 23716 33312
rect 23664 33269 23673 33303
rect 23673 33269 23707 33303
rect 23707 33269 23716 33303
rect 23664 33260 23716 33269
rect 25320 33260 25372 33312
rect 25688 33260 25740 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 6920 33056 6972 33108
rect 10784 33056 10836 33108
rect 12348 33056 12400 33108
rect 14464 33099 14516 33108
rect 14464 33065 14473 33099
rect 14473 33065 14507 33099
rect 14507 33065 14516 33099
rect 14464 33056 14516 33065
rect 16764 33056 16816 33108
rect 17500 33099 17552 33108
rect 17500 33065 17509 33099
rect 17509 33065 17543 33099
rect 17543 33065 17552 33099
rect 17500 33056 17552 33065
rect 19340 33056 19392 33108
rect 22192 33056 22244 33108
rect 23756 33099 23808 33108
rect 23756 33065 23765 33099
rect 23765 33065 23799 33099
rect 23799 33065 23808 33099
rect 23756 33056 23808 33065
rect 6736 32988 6788 33040
rect 10692 32988 10744 33040
rect 16488 32988 16540 33040
rect 6828 32920 6880 32972
rect 9864 32920 9916 32972
rect 9956 32920 10008 32972
rect 11888 32963 11940 32972
rect 11888 32929 11897 32963
rect 11897 32929 11931 32963
rect 11931 32929 11940 32963
rect 11888 32920 11940 32929
rect 13820 32963 13872 32972
rect 13820 32929 13829 32963
rect 13829 32929 13863 32963
rect 13863 32929 13872 32963
rect 13820 32920 13872 32929
rect 15016 32920 15068 32972
rect 18880 32920 18932 32972
rect 5448 32895 5500 32904
rect 5448 32861 5457 32895
rect 5457 32861 5491 32895
rect 5491 32861 5500 32895
rect 5448 32852 5500 32861
rect 5632 32852 5684 32904
rect 6460 32852 6512 32904
rect 9404 32852 9456 32904
rect 12348 32852 12400 32904
rect 13912 32852 13964 32904
rect 14096 32852 14148 32904
rect 14280 32895 14332 32904
rect 14280 32861 14289 32895
rect 14289 32861 14323 32895
rect 14323 32861 14332 32895
rect 14280 32852 14332 32861
rect 17684 32895 17736 32904
rect 17684 32861 17693 32895
rect 17693 32861 17727 32895
rect 17727 32861 17736 32895
rect 17684 32852 17736 32861
rect 7196 32784 7248 32836
rect 14372 32784 14424 32836
rect 16764 32784 16816 32836
rect 17776 32784 17828 32836
rect 19708 32988 19760 33040
rect 21180 32963 21232 32972
rect 21180 32929 21189 32963
rect 21189 32929 21223 32963
rect 21223 32929 21232 32963
rect 21180 32920 21232 32929
rect 23848 32988 23900 33040
rect 23296 32920 23348 32972
rect 23388 32920 23440 32972
rect 19708 32852 19760 32904
rect 19984 32895 20036 32904
rect 19984 32861 19993 32895
rect 19993 32861 20027 32895
rect 20027 32861 20036 32895
rect 19984 32852 20036 32861
rect 21916 32852 21968 32904
rect 22376 32852 22428 32904
rect 23664 32852 23716 32904
rect 25136 32895 25188 32904
rect 25136 32861 25145 32895
rect 25145 32861 25179 32895
rect 25179 32861 25188 32895
rect 25136 32852 25188 32861
rect 25780 32895 25832 32904
rect 25780 32861 25789 32895
rect 25789 32861 25823 32895
rect 25823 32861 25832 32895
rect 25780 32852 25832 32861
rect 12164 32759 12216 32768
rect 12164 32725 12173 32759
rect 12173 32725 12207 32759
rect 12207 32725 12216 32759
rect 12164 32716 12216 32725
rect 15752 32759 15804 32768
rect 15752 32725 15761 32759
rect 15761 32725 15795 32759
rect 15795 32725 15804 32759
rect 15752 32716 15804 32725
rect 18604 32716 18656 32768
rect 20168 32716 20220 32768
rect 23664 32716 23716 32768
rect 24676 32716 24728 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 6460 32555 6512 32564
rect 6460 32521 6469 32555
rect 6469 32521 6503 32555
rect 6503 32521 6512 32555
rect 6460 32512 6512 32521
rect 10600 32512 10652 32564
rect 11704 32512 11756 32564
rect 12072 32512 12124 32564
rect 5540 32419 5592 32428
rect 5540 32385 5549 32419
rect 5549 32385 5583 32419
rect 5583 32385 5592 32419
rect 5540 32376 5592 32385
rect 5724 32419 5776 32428
rect 5724 32385 5753 32419
rect 5753 32385 5776 32419
rect 5724 32376 5776 32385
rect 6644 32376 6696 32428
rect 7932 32376 7984 32428
rect 10140 32444 10192 32496
rect 10784 32444 10836 32496
rect 10876 32419 10928 32428
rect 10876 32385 10885 32419
rect 10885 32385 10919 32419
rect 10919 32385 10928 32419
rect 10876 32376 10928 32385
rect 12532 32512 12584 32564
rect 15752 32512 15804 32564
rect 16396 32512 16448 32564
rect 17684 32512 17736 32564
rect 19616 32512 19668 32564
rect 21916 32555 21968 32564
rect 21916 32521 21925 32555
rect 21925 32521 21959 32555
rect 21959 32521 21968 32555
rect 21916 32512 21968 32521
rect 23848 32555 23900 32564
rect 23848 32521 23857 32555
rect 23857 32521 23891 32555
rect 23891 32521 23900 32555
rect 23848 32512 23900 32521
rect 13820 32444 13872 32496
rect 17040 32444 17092 32496
rect 13084 32376 13136 32428
rect 15016 32419 15068 32428
rect 15016 32385 15025 32419
rect 15025 32385 15059 32419
rect 15059 32385 15068 32419
rect 15016 32376 15068 32385
rect 15292 32419 15344 32428
rect 15292 32385 15326 32419
rect 15326 32385 15344 32419
rect 15292 32376 15344 32385
rect 18880 32419 18932 32428
rect 18880 32385 18889 32419
rect 18889 32385 18923 32419
rect 18923 32385 18932 32419
rect 18880 32376 18932 32385
rect 19984 32376 20036 32428
rect 22376 32376 22428 32428
rect 23388 32444 23440 32496
rect 25136 32555 25188 32564
rect 25136 32521 25145 32555
rect 25145 32521 25179 32555
rect 25179 32521 25188 32555
rect 25136 32512 25188 32521
rect 848 32172 900 32224
rect 5632 32172 5684 32224
rect 7196 32172 7248 32224
rect 11060 32240 11112 32292
rect 14188 32240 14240 32292
rect 21916 32308 21968 32360
rect 23296 32376 23348 32428
rect 23664 32419 23716 32428
rect 23664 32385 23673 32419
rect 23673 32385 23707 32419
rect 23707 32385 23716 32419
rect 23664 32376 23716 32385
rect 24216 32376 24268 32428
rect 25688 32419 25740 32428
rect 23572 32351 23624 32360
rect 23572 32317 23581 32351
rect 23581 32317 23615 32351
rect 23615 32317 23624 32351
rect 23572 32308 23624 32317
rect 24676 32351 24728 32360
rect 24676 32317 24685 32351
rect 24685 32317 24719 32351
rect 24719 32317 24728 32351
rect 24676 32308 24728 32317
rect 19432 32240 19484 32292
rect 23848 32240 23900 32292
rect 25688 32385 25697 32419
rect 25697 32385 25731 32419
rect 25731 32385 25740 32419
rect 25688 32376 25740 32385
rect 27068 32419 27120 32428
rect 27068 32385 27077 32419
rect 27077 32385 27111 32419
rect 27111 32385 27120 32419
rect 27068 32376 27120 32385
rect 28264 32351 28316 32360
rect 28264 32317 28273 32351
rect 28273 32317 28307 32351
rect 28307 32317 28316 32351
rect 28264 32308 28316 32317
rect 12256 32172 12308 32224
rect 18788 32172 18840 32224
rect 22192 32172 22244 32224
rect 23112 32215 23164 32224
rect 23112 32181 23121 32215
rect 23121 32181 23155 32215
rect 23155 32181 23164 32215
rect 23112 32172 23164 32181
rect 25044 32172 25096 32224
rect 25136 32172 25188 32224
rect 25780 32172 25832 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 6000 31968 6052 32020
rect 7932 32011 7984 32020
rect 7932 31977 7941 32011
rect 7941 31977 7975 32011
rect 7975 31977 7984 32011
rect 7932 31968 7984 31977
rect 12716 32011 12768 32020
rect 12716 31977 12725 32011
rect 12725 31977 12759 32011
rect 12759 31977 12768 32011
rect 12716 31968 12768 31977
rect 15292 31968 15344 32020
rect 17040 31968 17092 32020
rect 18604 32011 18656 32020
rect 18604 31977 18613 32011
rect 18613 31977 18647 32011
rect 18647 31977 18656 32011
rect 18604 31968 18656 31977
rect 21088 31968 21140 32020
rect 21180 32011 21232 32020
rect 21180 31977 21189 32011
rect 21189 31977 21223 32011
rect 21223 31977 21232 32011
rect 21180 31968 21232 31977
rect 23756 31968 23808 32020
rect 7196 31764 7248 31816
rect 16396 31832 16448 31884
rect 19248 31832 19300 31884
rect 19708 31875 19760 31884
rect 19708 31841 19717 31875
rect 19717 31841 19751 31875
rect 19751 31841 19760 31875
rect 19708 31832 19760 31841
rect 22192 31832 22244 31884
rect 5632 31739 5684 31748
rect 5632 31705 5666 31739
rect 5666 31705 5684 31739
rect 5632 31696 5684 31705
rect 6644 31696 6696 31748
rect 8300 31807 8352 31816
rect 8300 31773 8309 31807
rect 8309 31773 8343 31807
rect 8343 31773 8352 31807
rect 8300 31764 8352 31773
rect 12164 31764 12216 31816
rect 12808 31807 12860 31816
rect 12808 31773 12817 31807
rect 12817 31773 12851 31807
rect 12851 31773 12860 31807
rect 12808 31764 12860 31773
rect 16488 31807 16540 31816
rect 16488 31773 16497 31807
rect 16497 31773 16531 31807
rect 16531 31773 16540 31807
rect 16488 31764 16540 31773
rect 18788 31807 18840 31816
rect 18788 31773 18797 31807
rect 18797 31773 18831 31807
rect 18831 31773 18840 31807
rect 18788 31764 18840 31773
rect 18880 31807 18932 31816
rect 18880 31773 18889 31807
rect 18889 31773 18923 31807
rect 18923 31773 18932 31807
rect 18880 31764 18932 31773
rect 18604 31739 18656 31748
rect 18604 31705 18613 31739
rect 18613 31705 18647 31739
rect 18647 31705 18656 31739
rect 18604 31696 18656 31705
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 19616 31807 19668 31816
rect 19616 31773 19625 31807
rect 19625 31773 19659 31807
rect 19659 31773 19668 31807
rect 19616 31764 19668 31773
rect 20812 31696 20864 31748
rect 21088 31764 21140 31816
rect 21456 31807 21508 31816
rect 21456 31773 21465 31807
rect 21465 31773 21499 31807
rect 21499 31773 21508 31807
rect 21456 31764 21508 31773
rect 21180 31696 21232 31748
rect 22008 31807 22060 31816
rect 22008 31773 22017 31807
rect 22017 31773 22051 31807
rect 22051 31773 22060 31807
rect 22008 31764 22060 31773
rect 22100 31807 22152 31816
rect 22100 31773 22109 31807
rect 22109 31773 22143 31807
rect 22143 31773 22152 31807
rect 22100 31764 22152 31773
rect 22744 31807 22796 31816
rect 22744 31773 22753 31807
rect 22753 31773 22787 31807
rect 22787 31773 22796 31807
rect 22744 31764 22796 31773
rect 23572 31764 23624 31816
rect 24584 31764 24636 31816
rect 28448 31807 28500 31816
rect 28448 31773 28457 31807
rect 28457 31773 28491 31807
rect 28491 31773 28500 31807
rect 28448 31764 28500 31773
rect 22100 31628 22152 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 8300 31424 8352 31476
rect 22744 31424 22796 31476
rect 20812 31356 20864 31408
rect 21916 31399 21968 31408
rect 21916 31365 21925 31399
rect 21925 31365 21959 31399
rect 21959 31365 21968 31399
rect 21916 31356 21968 31365
rect 22100 31399 22152 31408
rect 22100 31365 22109 31399
rect 22109 31365 22143 31399
rect 22143 31365 22152 31399
rect 22100 31356 22152 31365
rect 5908 31288 5960 31340
rect 6644 31331 6696 31340
rect 6644 31297 6653 31331
rect 6653 31297 6687 31331
rect 6687 31297 6696 31331
rect 6644 31288 6696 31297
rect 6828 31288 6880 31340
rect 21180 31331 21232 31340
rect 21180 31297 21189 31331
rect 21189 31297 21223 31331
rect 21223 31297 21232 31331
rect 21180 31288 21232 31297
rect 21456 31220 21508 31272
rect 22008 31220 22060 31272
rect 21548 31195 21600 31204
rect 21548 31161 21557 31195
rect 21557 31161 21591 31195
rect 21591 31161 21600 31195
rect 21548 31152 21600 31161
rect 6828 31127 6880 31136
rect 6828 31093 6837 31127
rect 6837 31093 6871 31127
rect 6871 31093 6880 31127
rect 6828 31084 6880 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 6736 30880 6788 30932
rect 18604 30923 18656 30932
rect 18604 30889 18613 30923
rect 18613 30889 18647 30923
rect 18647 30889 18656 30923
rect 18604 30880 18656 30889
rect 6828 30676 6880 30728
rect 7196 30676 7248 30728
rect 19616 30744 19668 30796
rect 17684 30608 17736 30660
rect 19248 30676 19300 30728
rect 6644 30540 6696 30592
rect 8484 30540 8536 30592
rect 17776 30540 17828 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 18604 30268 18656 30320
rect 24216 30311 24268 30320
rect 24216 30277 24225 30311
rect 24225 30277 24259 30311
rect 24259 30277 24268 30311
rect 24216 30268 24268 30277
rect 1308 30200 1360 30252
rect 9036 30132 9088 30184
rect 17684 30200 17736 30252
rect 19616 30200 19668 30252
rect 23756 30243 23808 30252
rect 23756 30209 23765 30243
rect 23765 30209 23799 30243
rect 23799 30209 23808 30243
rect 23756 30200 23808 30209
rect 23848 30243 23900 30252
rect 23848 30209 23857 30243
rect 23857 30209 23891 30243
rect 23891 30209 23900 30243
rect 23848 30200 23900 30209
rect 24124 30200 24176 30252
rect 19340 30132 19392 30184
rect 17316 30064 17368 30116
rect 17776 30064 17828 30116
rect 20628 30064 20680 30116
rect 1676 30039 1728 30048
rect 1676 30005 1685 30039
rect 1685 30005 1719 30039
rect 1719 30005 1728 30039
rect 1676 29996 1728 30005
rect 8484 29996 8536 30048
rect 9404 30039 9456 30048
rect 9404 30005 9413 30039
rect 9413 30005 9447 30039
rect 9447 30005 9456 30039
rect 9404 29996 9456 30005
rect 17500 30039 17552 30048
rect 17500 30005 17509 30039
rect 17509 30005 17543 30039
rect 17543 30005 17552 30039
rect 17500 29996 17552 30005
rect 18604 30039 18656 30048
rect 18604 30005 18613 30039
rect 18613 30005 18647 30039
rect 18647 30005 18656 30039
rect 18604 29996 18656 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 15108 29792 15160 29844
rect 17316 29792 17368 29844
rect 18788 29792 18840 29844
rect 19340 29835 19392 29844
rect 19340 29801 19349 29835
rect 19349 29801 19383 29835
rect 19383 29801 19392 29835
rect 19340 29792 19392 29801
rect 24584 29835 24636 29844
rect 24584 29801 24593 29835
rect 24593 29801 24627 29835
rect 24627 29801 24636 29835
rect 24584 29792 24636 29801
rect 9036 29767 9088 29776
rect 9036 29733 9045 29767
rect 9045 29733 9079 29767
rect 9079 29733 9088 29767
rect 9036 29724 9088 29733
rect 10508 29656 10560 29708
rect 17592 29699 17644 29708
rect 17592 29665 17601 29699
rect 17601 29665 17635 29699
rect 17635 29665 17644 29699
rect 17592 29656 17644 29665
rect 18604 29656 18656 29708
rect 19892 29699 19944 29708
rect 19892 29665 19901 29699
rect 19901 29665 19935 29699
rect 19935 29665 19944 29699
rect 19892 29656 19944 29665
rect 21916 29656 21968 29708
rect 848 29588 900 29640
rect 8484 29631 8536 29640
rect 8484 29597 8493 29631
rect 8493 29597 8527 29631
rect 8527 29597 8536 29631
rect 8484 29588 8536 29597
rect 10324 29588 10376 29640
rect 17500 29588 17552 29640
rect 24952 29520 25004 29572
rect 19432 29452 19484 29504
rect 24124 29495 24176 29504
rect 24124 29461 24133 29495
rect 24133 29461 24167 29495
rect 24167 29461 24176 29495
rect 24124 29452 24176 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 9772 29248 9824 29300
rect 10508 29248 10560 29300
rect 19616 29248 19668 29300
rect 8300 29180 8352 29232
rect 1676 29112 1728 29164
rect 8484 29112 8536 29164
rect 10876 29180 10928 29232
rect 12900 29180 12952 29232
rect 13544 29180 13596 29232
rect 12992 29155 13044 29164
rect 12992 29121 13001 29155
rect 13001 29121 13035 29155
rect 13035 29121 13044 29155
rect 12992 29112 13044 29121
rect 13636 29112 13688 29164
rect 13820 29112 13872 29164
rect 15108 29155 15160 29164
rect 15108 29121 15117 29155
rect 15117 29121 15151 29155
rect 15151 29121 15160 29155
rect 15108 29112 15160 29121
rect 15292 29155 15344 29164
rect 15292 29121 15301 29155
rect 15301 29121 15335 29155
rect 15335 29121 15344 29155
rect 15292 29112 15344 29121
rect 16396 29112 16448 29164
rect 18144 29180 18196 29232
rect 16764 29155 16816 29164
rect 16764 29121 16773 29155
rect 16773 29121 16807 29155
rect 16807 29121 16816 29155
rect 16764 29112 16816 29121
rect 16948 29155 17000 29164
rect 16948 29121 16957 29155
rect 16957 29121 16991 29155
rect 16991 29121 17000 29155
rect 16948 29112 17000 29121
rect 4804 28976 4856 29028
rect 10048 28976 10100 29028
rect 9864 28908 9916 28960
rect 10324 28908 10376 28960
rect 10968 28908 11020 28960
rect 11336 29044 11388 29096
rect 15200 29087 15252 29096
rect 15200 29053 15209 29087
rect 15209 29053 15243 29087
rect 15243 29053 15252 29087
rect 15200 29044 15252 29053
rect 17960 29044 18012 29096
rect 21916 29180 21968 29232
rect 24952 29248 25004 29300
rect 27068 29248 27120 29300
rect 24124 29180 24176 29232
rect 18788 29112 18840 29164
rect 19432 29044 19484 29096
rect 23664 29087 23716 29096
rect 23664 29053 23673 29087
rect 23673 29053 23707 29087
rect 23707 29053 23716 29087
rect 23664 29044 23716 29053
rect 25320 29155 25372 29164
rect 25320 29121 25329 29155
rect 25329 29121 25363 29155
rect 25363 29121 25372 29155
rect 25320 29112 25372 29121
rect 26056 29112 26108 29164
rect 14372 28976 14424 29028
rect 14740 28976 14792 29028
rect 16764 28976 16816 29028
rect 11428 28908 11480 28960
rect 17040 28908 17092 28960
rect 19892 28976 19944 29028
rect 23848 28976 23900 29028
rect 19524 28908 19576 28960
rect 24032 28951 24084 28960
rect 24032 28917 24041 28951
rect 24041 28917 24075 28951
rect 24075 28917 24084 28951
rect 24032 28908 24084 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 10140 28704 10192 28756
rect 11336 28704 11388 28756
rect 11060 28636 11112 28688
rect 12992 28704 13044 28756
rect 15292 28704 15344 28756
rect 16856 28704 16908 28756
rect 17500 28704 17552 28756
rect 26056 28747 26108 28756
rect 26056 28713 26065 28747
rect 26065 28713 26099 28747
rect 26099 28713 26108 28747
rect 26056 28704 26108 28713
rect 17684 28679 17736 28688
rect 17684 28645 17693 28679
rect 17693 28645 17727 28679
rect 17727 28645 17736 28679
rect 17684 28636 17736 28645
rect 9404 28568 9456 28620
rect 4804 28475 4856 28484
rect 4804 28441 4838 28475
rect 4838 28441 4856 28475
rect 4804 28432 4856 28441
rect 7196 28432 7248 28484
rect 8300 28500 8352 28552
rect 9772 28568 9824 28620
rect 9864 28611 9916 28620
rect 9864 28577 9873 28611
rect 9873 28577 9907 28611
rect 9907 28577 9916 28611
rect 9864 28568 9916 28577
rect 13084 28568 13136 28620
rect 21548 28568 21600 28620
rect 8668 28475 8720 28484
rect 8668 28441 8677 28475
rect 8677 28441 8711 28475
rect 8711 28441 8720 28475
rect 8668 28432 8720 28441
rect 9128 28432 9180 28484
rect 10048 28432 10100 28484
rect 14096 28500 14148 28552
rect 12348 28475 12400 28484
rect 12348 28441 12382 28475
rect 12382 28441 12400 28475
rect 12348 28432 12400 28441
rect 13820 28432 13872 28484
rect 6828 28364 6880 28416
rect 7472 28364 7524 28416
rect 8208 28407 8260 28416
rect 8208 28373 8217 28407
rect 8217 28373 8251 28407
rect 8251 28373 8260 28407
rect 8208 28364 8260 28373
rect 8484 28364 8536 28416
rect 9312 28407 9364 28416
rect 9312 28373 9321 28407
rect 9321 28373 9355 28407
rect 9355 28373 9364 28407
rect 9312 28364 9364 28373
rect 9404 28407 9456 28416
rect 9404 28373 9413 28407
rect 9413 28373 9447 28407
rect 9447 28373 9456 28407
rect 9404 28364 9456 28373
rect 9956 28364 10008 28416
rect 13636 28364 13688 28416
rect 14648 28543 14700 28552
rect 14648 28509 14657 28543
rect 14657 28509 14691 28543
rect 14691 28509 14700 28543
rect 14648 28500 14700 28509
rect 16580 28543 16632 28552
rect 16580 28509 16589 28543
rect 16589 28509 16623 28543
rect 16623 28509 16632 28543
rect 16580 28500 16632 28509
rect 16672 28500 16724 28552
rect 17132 28543 17184 28552
rect 17132 28509 17141 28543
rect 17141 28509 17175 28543
rect 17175 28509 17184 28543
rect 17132 28500 17184 28509
rect 17776 28500 17828 28552
rect 19524 28543 19576 28552
rect 19524 28509 19533 28543
rect 19533 28509 19567 28543
rect 19567 28509 19576 28543
rect 19524 28500 19576 28509
rect 19892 28500 19944 28552
rect 23848 28568 23900 28620
rect 24860 28568 24912 28620
rect 23204 28500 23256 28552
rect 23664 28500 23716 28552
rect 24492 28500 24544 28552
rect 17684 28432 17736 28484
rect 24584 28432 24636 28484
rect 19432 28407 19484 28416
rect 19432 28373 19441 28407
rect 19441 28373 19475 28407
rect 19475 28373 19484 28407
rect 19432 28364 19484 28373
rect 20904 28407 20956 28416
rect 20904 28373 20913 28407
rect 20913 28373 20947 28407
rect 20947 28373 20956 28407
rect 20904 28364 20956 28373
rect 21548 28407 21600 28416
rect 21548 28373 21557 28407
rect 21557 28373 21591 28407
rect 21591 28373 21600 28407
rect 21548 28364 21600 28373
rect 23480 28364 23532 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 8484 28160 8536 28212
rect 10048 28203 10100 28212
rect 10048 28169 10057 28203
rect 10057 28169 10091 28203
rect 10091 28169 10100 28203
rect 10048 28160 10100 28169
rect 10508 28160 10560 28212
rect 10876 28203 10928 28212
rect 10876 28169 10885 28203
rect 10885 28169 10919 28203
rect 10919 28169 10928 28203
rect 10876 28160 10928 28169
rect 13084 28160 13136 28212
rect 15384 28203 15436 28212
rect 15384 28169 15393 28203
rect 15393 28169 15427 28203
rect 15427 28169 15436 28203
rect 15384 28160 15436 28169
rect 6828 28067 6880 28076
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 14188 28092 14240 28144
rect 7472 28067 7524 28076
rect 7472 28033 7506 28067
rect 7506 28033 7524 28067
rect 7472 28024 7524 28033
rect 9956 28067 10008 28076
rect 9956 28033 9965 28067
rect 9965 28033 9999 28067
rect 9999 28033 10008 28067
rect 9956 28024 10008 28033
rect 10140 28024 10192 28076
rect 11060 28067 11112 28076
rect 11060 28033 11069 28067
rect 11069 28033 11103 28067
rect 11103 28033 11112 28067
rect 11060 28024 11112 28033
rect 112 27888 164 27940
rect 7196 27999 7248 28008
rect 7196 27965 7205 27999
rect 7205 27965 7239 27999
rect 7239 27965 7248 27999
rect 7196 27956 7248 27965
rect 8668 27888 8720 27940
rect 10968 27956 11020 28008
rect 12164 28024 12216 28076
rect 12716 28024 12768 28076
rect 11428 27956 11480 28008
rect 13360 27999 13412 28008
rect 13360 27965 13369 27999
rect 13369 27965 13403 27999
rect 13403 27965 13412 27999
rect 13360 27956 13412 27965
rect 10508 27888 10560 27940
rect 6736 27820 6788 27872
rect 8852 27863 8904 27872
rect 8852 27829 8861 27863
rect 8861 27829 8895 27863
rect 8895 27829 8904 27863
rect 8852 27820 8904 27829
rect 10876 27820 10928 27872
rect 14004 27888 14056 27940
rect 16948 28160 17000 28212
rect 22100 28203 22152 28212
rect 22100 28169 22109 28203
rect 22109 28169 22143 28203
rect 22143 28169 22152 28203
rect 22100 28160 22152 28169
rect 24032 28203 24084 28212
rect 24032 28169 24041 28203
rect 24041 28169 24075 28203
rect 24075 28169 24084 28203
rect 24032 28160 24084 28169
rect 24492 28203 24544 28212
rect 24492 28169 24501 28203
rect 24501 28169 24535 28203
rect 24535 28169 24544 28203
rect 24492 28160 24544 28169
rect 24584 28160 24636 28212
rect 16672 28024 16724 28076
rect 17684 28024 17736 28076
rect 17960 28067 18012 28076
rect 17960 28033 17969 28067
rect 17969 28033 18003 28067
rect 18003 28033 18012 28067
rect 17960 28024 18012 28033
rect 20904 28067 20956 28076
rect 20904 28033 20913 28067
rect 20913 28033 20947 28067
rect 20947 28033 20956 28067
rect 20904 28024 20956 28033
rect 17408 27956 17460 28008
rect 20628 27999 20680 28008
rect 20628 27965 20637 27999
rect 20637 27965 20671 27999
rect 20671 27965 20680 27999
rect 22192 28024 22244 28076
rect 23112 28024 23164 28076
rect 23480 28067 23532 28076
rect 23480 28033 23489 28067
rect 23489 28033 23523 28067
rect 23523 28033 23532 28067
rect 23480 28024 23532 28033
rect 24032 28024 24084 28076
rect 24952 28067 25004 28076
rect 24952 28033 24961 28067
rect 24961 28033 24995 28067
rect 24995 28033 25004 28067
rect 24952 28024 25004 28033
rect 20628 27956 20680 27965
rect 23848 27999 23900 28008
rect 23848 27965 23857 27999
rect 23857 27965 23891 27999
rect 23891 27965 23900 27999
rect 23848 27956 23900 27965
rect 17224 27888 17276 27940
rect 12348 27820 12400 27872
rect 20904 27863 20956 27872
rect 20904 27829 20913 27863
rect 20913 27829 20947 27863
rect 20947 27829 20956 27863
rect 20904 27820 20956 27829
rect 21548 27820 21600 27872
rect 22008 27820 22060 27872
rect 23480 27863 23532 27872
rect 23480 27829 23489 27863
rect 23489 27829 23523 27863
rect 23523 27829 23532 27863
rect 23480 27820 23532 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 9312 27616 9364 27668
rect 12164 27659 12216 27668
rect 12164 27625 12173 27659
rect 12173 27625 12207 27659
rect 12207 27625 12216 27659
rect 12164 27616 12216 27625
rect 12716 27659 12768 27668
rect 12716 27625 12725 27659
rect 12725 27625 12759 27659
rect 12759 27625 12768 27659
rect 12716 27616 12768 27625
rect 14188 27659 14240 27668
rect 14188 27625 14197 27659
rect 14197 27625 14231 27659
rect 14231 27625 14240 27659
rect 14188 27616 14240 27625
rect 8300 27548 8352 27600
rect 8392 27523 8444 27532
rect 8392 27489 8401 27523
rect 8401 27489 8435 27523
rect 8435 27489 8444 27523
rect 8392 27480 8444 27489
rect 9404 27480 9456 27532
rect 13084 27480 13136 27532
rect 14096 27480 14148 27532
rect 17592 27616 17644 27668
rect 17684 27659 17736 27668
rect 17684 27625 17693 27659
rect 17693 27625 17727 27659
rect 17727 27625 17736 27659
rect 17684 27616 17736 27625
rect 22192 27659 22244 27668
rect 22192 27625 22201 27659
rect 22201 27625 22235 27659
rect 22235 27625 22244 27659
rect 22192 27616 22244 27625
rect 24952 27616 25004 27668
rect 16580 27548 16632 27600
rect 17500 27591 17552 27600
rect 17500 27557 17509 27591
rect 17509 27557 17543 27591
rect 17543 27557 17552 27591
rect 17500 27548 17552 27557
rect 16764 27480 16816 27532
rect 17040 27523 17092 27532
rect 17040 27489 17049 27523
rect 17049 27489 17083 27523
rect 17083 27489 17092 27523
rect 17040 27480 17092 27489
rect 7196 27412 7248 27464
rect 8208 27455 8260 27464
rect 8208 27421 8217 27455
rect 8217 27421 8251 27455
rect 8251 27421 8260 27455
rect 8208 27412 8260 27421
rect 9128 27412 9180 27464
rect 10048 27455 10100 27464
rect 10048 27421 10057 27455
rect 10057 27421 10091 27455
rect 10091 27421 10100 27455
rect 10048 27412 10100 27421
rect 11060 27412 11112 27464
rect 16856 27455 16908 27464
rect 16856 27421 16865 27455
rect 16865 27421 16899 27455
rect 16899 27421 16908 27455
rect 16856 27412 16908 27421
rect 17132 27412 17184 27464
rect 18144 27455 18196 27464
rect 18144 27421 18153 27455
rect 18153 27421 18187 27455
rect 18187 27421 18196 27455
rect 18144 27412 18196 27421
rect 21456 27412 21508 27464
rect 23480 27412 23532 27464
rect 28448 27455 28500 27464
rect 28448 27421 28457 27455
rect 28457 27421 28491 27455
rect 28491 27421 28500 27455
rect 28448 27412 28500 27421
rect 6736 27387 6788 27396
rect 6736 27353 6770 27387
rect 6770 27353 6788 27387
rect 6736 27344 6788 27353
rect 15200 27344 15252 27396
rect 10692 27276 10744 27328
rect 16672 27344 16724 27396
rect 17868 27387 17920 27396
rect 17868 27353 17877 27387
rect 17877 27353 17911 27387
rect 17911 27353 17920 27387
rect 17868 27344 17920 27353
rect 20904 27344 20956 27396
rect 16764 27276 16816 27328
rect 17132 27276 17184 27328
rect 17776 27276 17828 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 8392 27115 8444 27124
rect 8392 27081 8401 27115
rect 8401 27081 8435 27115
rect 8435 27081 8444 27115
rect 8392 27072 8444 27081
rect 10048 27115 10100 27124
rect 10048 27081 10057 27115
rect 10057 27081 10091 27115
rect 10091 27081 10100 27115
rect 10048 27072 10100 27081
rect 11060 27115 11112 27124
rect 11060 27081 11069 27115
rect 11069 27081 11103 27115
rect 11103 27081 11112 27115
rect 11060 27072 11112 27081
rect 12348 27072 12400 27124
rect 7196 27004 7248 27056
rect 8116 26936 8168 26988
rect 9864 27004 9916 27056
rect 10692 27047 10744 27056
rect 10692 27013 10701 27047
rect 10701 27013 10735 27047
rect 10735 27013 10744 27047
rect 10692 27004 10744 27013
rect 11428 27004 11480 27056
rect 12992 27072 13044 27124
rect 16672 27072 16724 27124
rect 17408 27115 17460 27124
rect 17408 27081 17417 27115
rect 17417 27081 17451 27115
rect 17451 27081 17460 27115
rect 17408 27072 17460 27081
rect 22376 27072 22428 27124
rect 8944 26979 8996 26988
rect 8944 26945 8978 26979
rect 8978 26945 8996 26979
rect 8944 26936 8996 26945
rect 10508 26979 10560 26988
rect 10508 26945 10517 26979
rect 10517 26945 10551 26979
rect 10551 26945 10560 26979
rect 10508 26936 10560 26945
rect 10876 26979 10928 26988
rect 10876 26945 10885 26979
rect 10885 26945 10919 26979
rect 10919 26945 10928 26979
rect 10876 26936 10928 26945
rect 12716 26936 12768 26988
rect 13084 26936 13136 26988
rect 13912 27004 13964 27056
rect 14648 27004 14700 27056
rect 13820 26979 13872 26988
rect 13820 26945 13829 26979
rect 13829 26945 13863 26979
rect 13863 26945 13872 26979
rect 13820 26936 13872 26945
rect 14004 26936 14056 26988
rect 14740 26979 14792 26988
rect 14740 26945 14749 26979
rect 14749 26945 14783 26979
rect 14783 26945 14792 26979
rect 14740 26936 14792 26945
rect 20260 27004 20312 27056
rect 24032 27072 24084 27124
rect 25136 27115 25188 27124
rect 25136 27081 25145 27115
rect 25145 27081 25179 27115
rect 25179 27081 25188 27115
rect 25136 27072 25188 27081
rect 16764 26979 16816 26988
rect 16764 26945 16773 26979
rect 16773 26945 16807 26979
rect 16807 26945 16816 26979
rect 16764 26936 16816 26945
rect 17960 26936 18012 26988
rect 14372 26868 14424 26920
rect 16856 26868 16908 26920
rect 17684 26868 17736 26920
rect 18604 26979 18656 26988
rect 18604 26945 18613 26979
rect 18613 26945 18647 26979
rect 18647 26945 18656 26979
rect 18604 26936 18656 26945
rect 20628 26936 20680 26988
rect 22008 26979 22060 26988
rect 22008 26945 22018 26979
rect 22018 26945 22052 26979
rect 22052 26945 22060 26979
rect 22008 26936 22060 26945
rect 22284 26868 22336 26920
rect 17040 26800 17092 26852
rect 23020 26979 23072 26988
rect 23020 26945 23029 26979
rect 23029 26945 23063 26979
rect 23063 26945 23072 26979
rect 23020 26936 23072 26945
rect 23940 26979 23992 26988
rect 23940 26945 23949 26979
rect 23949 26945 23983 26979
rect 23983 26945 23992 26979
rect 23940 26936 23992 26945
rect 24032 26979 24084 26988
rect 24032 26945 24041 26979
rect 24041 26945 24075 26979
rect 24075 26945 24084 26979
rect 24032 26936 24084 26945
rect 25228 26979 25280 26988
rect 25228 26945 25237 26979
rect 25237 26945 25271 26979
rect 25271 26945 25280 26979
rect 25228 26936 25280 26945
rect 25228 26800 25280 26852
rect 13636 26775 13688 26784
rect 13636 26741 13645 26775
rect 13645 26741 13679 26775
rect 13679 26741 13688 26775
rect 13636 26732 13688 26741
rect 19892 26732 19944 26784
rect 24860 26775 24912 26784
rect 24860 26741 24869 26775
rect 24869 26741 24903 26775
rect 24903 26741 24912 26775
rect 24860 26732 24912 26741
rect 24952 26775 25004 26784
rect 24952 26741 24961 26775
rect 24961 26741 24995 26775
rect 24995 26741 25004 26775
rect 24952 26732 25004 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 8116 26571 8168 26580
rect 8116 26537 8125 26571
rect 8125 26537 8159 26571
rect 8159 26537 8168 26571
rect 8116 26528 8168 26537
rect 13820 26571 13872 26580
rect 13820 26537 13829 26571
rect 13829 26537 13863 26571
rect 13863 26537 13872 26571
rect 13820 26528 13872 26537
rect 17684 26571 17736 26580
rect 17684 26537 17693 26571
rect 17693 26537 17727 26571
rect 17727 26537 17736 26571
rect 17684 26528 17736 26537
rect 17960 26571 18012 26580
rect 17960 26537 17969 26571
rect 17969 26537 18003 26571
rect 18003 26537 18012 26571
rect 17960 26528 18012 26537
rect 20628 26571 20680 26580
rect 20628 26537 20637 26571
rect 20637 26537 20671 26571
rect 20671 26537 20680 26571
rect 20628 26528 20680 26537
rect 23020 26528 23072 26580
rect 8852 26392 8904 26444
rect 9404 26392 9456 26444
rect 19156 26392 19208 26444
rect 20168 26435 20220 26444
rect 20168 26401 20177 26435
rect 20177 26401 20211 26435
rect 20211 26401 20220 26435
rect 20168 26392 20220 26401
rect 20260 26435 20312 26444
rect 20260 26401 20269 26435
rect 20269 26401 20303 26435
rect 20303 26401 20312 26435
rect 20260 26392 20312 26401
rect 8300 26367 8352 26376
rect 8300 26333 8309 26367
rect 8309 26333 8343 26367
rect 8343 26333 8352 26367
rect 8300 26324 8352 26333
rect 12256 26324 12308 26376
rect 17132 26367 17184 26376
rect 17132 26333 17141 26367
rect 17141 26333 17175 26367
rect 17175 26333 17184 26367
rect 17132 26324 17184 26333
rect 18144 26367 18196 26376
rect 12716 26299 12768 26308
rect 12716 26265 12750 26299
rect 12750 26265 12768 26299
rect 12716 26256 12768 26265
rect 17040 26256 17092 26308
rect 18144 26333 18153 26367
rect 18153 26333 18187 26367
rect 18187 26333 18196 26367
rect 18144 26324 18196 26333
rect 17868 26256 17920 26308
rect 19432 26324 19484 26376
rect 19892 26367 19944 26376
rect 19892 26333 19901 26367
rect 19901 26333 19935 26367
rect 19935 26333 19944 26367
rect 19892 26324 19944 26333
rect 22008 26324 22060 26376
rect 22376 26324 22428 26376
rect 21180 26256 21232 26308
rect 22284 26299 22336 26308
rect 22284 26265 22293 26299
rect 22293 26265 22327 26299
rect 22327 26265 22336 26299
rect 22284 26256 22336 26265
rect 22836 26256 22888 26308
rect 9312 26188 9364 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 8944 25984 8996 26036
rect 12716 26027 12768 26036
rect 12716 25993 12725 26027
rect 12725 25993 12759 26027
rect 12759 25993 12768 26027
rect 12716 25984 12768 25993
rect 13360 26027 13412 26036
rect 8300 25644 8352 25696
rect 9312 25891 9364 25900
rect 9312 25857 9321 25891
rect 9321 25857 9355 25891
rect 9355 25857 9364 25891
rect 9312 25848 9364 25857
rect 13360 25993 13369 26027
rect 13369 25993 13403 26027
rect 13403 25993 13412 26027
rect 13360 25984 13412 25993
rect 18604 25984 18656 26036
rect 20996 25984 21048 26036
rect 21180 25984 21232 26036
rect 20168 25916 20220 25968
rect 9772 25687 9824 25696
rect 9772 25653 9781 25687
rect 9781 25653 9815 25687
rect 9815 25653 9824 25687
rect 19156 25891 19208 25900
rect 19156 25857 19165 25891
rect 19165 25857 19199 25891
rect 19199 25857 19208 25891
rect 19156 25848 19208 25857
rect 19432 25848 19484 25900
rect 13912 25823 13964 25832
rect 13912 25789 13921 25823
rect 13921 25789 13955 25823
rect 13955 25789 13964 25823
rect 13912 25780 13964 25789
rect 18604 25780 18656 25832
rect 25780 25823 25832 25832
rect 25780 25789 25789 25823
rect 25789 25789 25823 25823
rect 25823 25789 25832 25823
rect 25780 25780 25832 25789
rect 9772 25644 9824 25653
rect 24952 25644 25004 25696
rect 25228 25687 25280 25696
rect 25228 25653 25237 25687
rect 25237 25653 25271 25687
rect 25271 25653 25280 25687
rect 25228 25644 25280 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 21180 25440 21232 25492
rect 19800 25279 19852 25288
rect 19800 25245 19809 25279
rect 19809 25245 19843 25279
rect 19843 25245 19852 25279
rect 19800 25236 19852 25245
rect 20536 25236 20588 25288
rect 20904 25211 20956 25220
rect 20904 25177 20913 25211
rect 20913 25177 20947 25211
rect 20947 25177 20956 25211
rect 20904 25168 20956 25177
rect 19524 25100 19576 25152
rect 20720 25100 20772 25152
rect 21272 25143 21324 25152
rect 21272 25109 21281 25143
rect 21281 25109 21315 25143
rect 21315 25109 21324 25143
rect 21272 25100 21324 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 18052 24871 18104 24880
rect 18052 24837 18061 24871
rect 18061 24837 18095 24871
rect 18095 24837 18104 24871
rect 18052 24828 18104 24837
rect 12256 24760 12308 24812
rect 12440 24803 12492 24812
rect 12440 24769 12474 24803
rect 12474 24769 12492 24803
rect 12440 24760 12492 24769
rect 18236 24760 18288 24812
rect 19524 24803 19576 24812
rect 19524 24769 19533 24803
rect 19533 24769 19567 24803
rect 19567 24769 19576 24803
rect 19524 24760 19576 24769
rect 21180 24828 21232 24880
rect 23388 24871 23440 24880
rect 21088 24760 21140 24812
rect 22100 24803 22152 24812
rect 22100 24769 22109 24803
rect 22109 24769 22143 24803
rect 22143 24769 22152 24803
rect 22100 24760 22152 24769
rect 23388 24837 23397 24871
rect 23397 24837 23431 24871
rect 23431 24837 23440 24871
rect 23388 24828 23440 24837
rect 20076 24692 20128 24744
rect 20812 24692 20864 24744
rect 20996 24735 21048 24744
rect 20996 24701 21005 24735
rect 21005 24701 21039 24735
rect 21039 24701 21048 24735
rect 20996 24692 21048 24701
rect 23756 24760 23808 24812
rect 13912 24624 13964 24676
rect 18512 24624 18564 24676
rect 20720 24624 20772 24676
rect 21272 24624 21324 24676
rect 24124 24692 24176 24744
rect 17960 24556 18012 24608
rect 19432 24556 19484 24608
rect 19800 24556 19852 24608
rect 20628 24599 20680 24608
rect 20628 24565 20637 24599
rect 20637 24565 20671 24599
rect 20671 24565 20680 24599
rect 20628 24556 20680 24565
rect 21916 24599 21968 24608
rect 21916 24565 21925 24599
rect 21925 24565 21959 24599
rect 21959 24565 21968 24599
rect 21916 24556 21968 24565
rect 22652 24599 22704 24608
rect 22652 24565 22661 24599
rect 22661 24565 22695 24599
rect 22695 24565 22704 24599
rect 22652 24556 22704 24565
rect 23112 24556 23164 24608
rect 23572 24599 23624 24608
rect 23572 24565 23581 24599
rect 23581 24565 23615 24599
rect 23615 24565 23624 24599
rect 23572 24556 23624 24565
rect 24492 24556 24544 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 12440 24352 12492 24404
rect 20904 24352 20956 24404
rect 24676 24284 24728 24336
rect 17040 24259 17092 24268
rect 17040 24225 17049 24259
rect 17049 24225 17083 24259
rect 17083 24225 17092 24259
rect 17040 24216 17092 24225
rect 18236 24259 18288 24268
rect 848 24148 900 24200
rect 11060 24191 11112 24200
rect 11060 24157 11069 24191
rect 11069 24157 11103 24191
rect 11103 24157 11112 24191
rect 11060 24148 11112 24157
rect 11980 24148 12032 24200
rect 12624 24191 12676 24200
rect 12624 24157 12633 24191
rect 12633 24157 12667 24191
rect 12667 24157 12676 24191
rect 12624 24148 12676 24157
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 17592 24148 17644 24200
rect 18236 24225 18245 24259
rect 18245 24225 18279 24259
rect 18279 24225 18288 24259
rect 18236 24216 18288 24225
rect 20628 24259 20680 24268
rect 20628 24225 20637 24259
rect 20637 24225 20671 24259
rect 20671 24225 20680 24259
rect 20628 24216 20680 24225
rect 22652 24216 22704 24268
rect 23572 24216 23624 24268
rect 18052 24148 18104 24200
rect 18144 24148 18196 24200
rect 19340 24191 19392 24200
rect 19340 24157 19349 24191
rect 19349 24157 19383 24191
rect 19383 24157 19392 24191
rect 19340 24148 19392 24157
rect 20260 24148 20312 24200
rect 23756 24191 23808 24200
rect 23756 24157 23765 24191
rect 23765 24157 23799 24191
rect 23799 24157 23808 24191
rect 23756 24148 23808 24157
rect 24492 24191 24544 24200
rect 24492 24157 24501 24191
rect 24501 24157 24535 24191
rect 24535 24157 24544 24191
rect 24492 24148 24544 24157
rect 10600 24012 10652 24064
rect 16304 24012 16356 24064
rect 21272 24080 21324 24132
rect 24308 24080 24360 24132
rect 17316 24055 17368 24064
rect 17316 24021 17325 24055
rect 17325 24021 17359 24055
rect 17359 24021 17368 24055
rect 17316 24012 17368 24021
rect 19524 24012 19576 24064
rect 21180 24055 21232 24064
rect 21180 24021 21189 24055
rect 21189 24021 21223 24055
rect 21223 24021 21232 24055
rect 21180 24012 21232 24021
rect 22652 24055 22704 24064
rect 22652 24021 22661 24055
rect 22661 24021 22695 24055
rect 22695 24021 22704 24055
rect 22652 24012 22704 24021
rect 23112 24012 23164 24064
rect 24952 24012 25004 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 11060 23808 11112 23860
rect 12072 23808 12124 23860
rect 17500 23808 17552 23860
rect 18144 23851 18196 23860
rect 18144 23817 18153 23851
rect 18153 23817 18187 23851
rect 18187 23817 18196 23851
rect 18144 23808 18196 23817
rect 20260 23808 20312 23860
rect 23572 23808 23624 23860
rect 25780 23808 25832 23860
rect 16304 23783 16356 23792
rect 8760 23672 8812 23724
rect 9772 23672 9824 23724
rect 8484 23604 8536 23656
rect 10600 23715 10652 23724
rect 10600 23681 10609 23715
rect 10609 23681 10643 23715
rect 10643 23681 10652 23715
rect 10600 23672 10652 23681
rect 11980 23672 12032 23724
rect 12716 23672 12768 23724
rect 14464 23672 14516 23724
rect 15752 23672 15804 23724
rect 16304 23749 16313 23783
rect 16313 23749 16347 23783
rect 16347 23749 16356 23783
rect 16304 23740 16356 23749
rect 17316 23740 17368 23792
rect 19524 23783 19576 23792
rect 19524 23749 19542 23783
rect 19542 23749 19576 23783
rect 19524 23740 19576 23749
rect 12164 23647 12216 23656
rect 12164 23613 12173 23647
rect 12173 23613 12207 23647
rect 12207 23613 12216 23647
rect 12164 23604 12216 23613
rect 14280 23604 14332 23656
rect 17592 23672 17644 23724
rect 21180 23715 21232 23724
rect 21180 23681 21198 23715
rect 21198 23681 21232 23715
rect 21180 23672 21232 23681
rect 21456 23715 21508 23724
rect 21456 23681 21465 23715
rect 21465 23681 21499 23715
rect 21499 23681 21508 23715
rect 21456 23672 21508 23681
rect 24492 23672 24544 23724
rect 16764 23647 16816 23656
rect 16764 23613 16773 23647
rect 16773 23613 16807 23647
rect 16807 23613 16816 23647
rect 16764 23604 16816 23613
rect 21916 23604 21968 23656
rect 22836 23647 22888 23656
rect 22836 23613 22845 23647
rect 22845 23613 22879 23647
rect 22879 23613 22888 23647
rect 22836 23604 22888 23613
rect 13544 23536 13596 23588
rect 848 23468 900 23520
rect 10324 23511 10376 23520
rect 10324 23477 10333 23511
rect 10333 23477 10367 23511
rect 10367 23477 10376 23511
rect 10324 23468 10376 23477
rect 10876 23468 10928 23520
rect 13268 23468 13320 23520
rect 13636 23511 13688 23520
rect 13636 23477 13645 23511
rect 13645 23477 13679 23511
rect 13679 23477 13688 23511
rect 13636 23468 13688 23477
rect 15660 23511 15712 23520
rect 15660 23477 15669 23511
rect 15669 23477 15703 23511
rect 15703 23477 15712 23511
rect 15660 23468 15712 23477
rect 18604 23468 18656 23520
rect 21732 23468 21784 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 6460 23060 6512 23112
rect 8484 23128 8536 23180
rect 12164 23264 12216 23316
rect 12624 23264 12676 23316
rect 12072 23196 12124 23248
rect 4620 22992 4672 23044
rect 9404 23060 9456 23112
rect 11796 23060 11848 23112
rect 12808 23196 12860 23248
rect 13544 23196 13596 23248
rect 13728 23128 13780 23180
rect 14004 23128 14056 23180
rect 16764 23264 16816 23316
rect 17040 23196 17092 23248
rect 20996 23264 21048 23316
rect 21088 23264 21140 23316
rect 22836 23307 22888 23316
rect 22836 23273 22845 23307
rect 22845 23273 22879 23307
rect 22879 23273 22888 23307
rect 22836 23264 22888 23273
rect 23388 23264 23440 23316
rect 24492 23307 24544 23316
rect 24492 23273 24501 23307
rect 24501 23273 24535 23307
rect 24535 23273 24544 23307
rect 24492 23264 24544 23273
rect 24584 23264 24636 23316
rect 21456 23171 21508 23180
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 12624 23060 12676 23069
rect 12716 23103 12768 23112
rect 12716 23069 12725 23103
rect 12725 23069 12759 23103
rect 12759 23069 12768 23103
rect 12716 23060 12768 23069
rect 13268 23103 13320 23112
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 10324 23035 10376 23044
rect 10324 23001 10342 23035
rect 10342 23001 10376 23035
rect 10324 22992 10376 23001
rect 12164 22992 12216 23044
rect 14464 23103 14516 23112
rect 14464 23069 14473 23103
rect 14473 23069 14507 23103
rect 14507 23069 14516 23103
rect 14464 23060 14516 23069
rect 14648 23103 14700 23112
rect 14648 23069 14657 23103
rect 14657 23069 14691 23103
rect 14691 23069 14700 23103
rect 14648 23060 14700 23069
rect 15660 23060 15712 23112
rect 18144 23060 18196 23112
rect 18696 23060 18748 23112
rect 21456 23137 21465 23171
rect 21465 23137 21499 23171
rect 21499 23137 21508 23171
rect 21456 23128 21508 23137
rect 23940 23128 23992 23180
rect 24952 23171 25004 23180
rect 24952 23137 24961 23171
rect 24961 23137 24995 23171
rect 24995 23137 25004 23171
rect 24952 23128 25004 23137
rect 20536 23060 20588 23112
rect 17960 23035 18012 23044
rect 17960 23001 17969 23035
rect 17969 23001 18003 23035
rect 18003 23001 18012 23035
rect 17960 22992 18012 23001
rect 19432 22992 19484 23044
rect 21272 23060 21324 23112
rect 21732 23103 21784 23112
rect 21732 23069 21766 23103
rect 21766 23069 21784 23103
rect 21732 23060 21784 23069
rect 24676 23103 24728 23112
rect 24676 23069 24685 23103
rect 24685 23069 24719 23103
rect 24719 23069 24728 23103
rect 24676 23060 24728 23069
rect 23388 22992 23440 23044
rect 8392 22967 8444 22976
rect 8392 22933 8401 22967
rect 8401 22933 8435 22967
rect 8435 22933 8444 22967
rect 8392 22924 8444 22933
rect 9772 22924 9824 22976
rect 11612 22967 11664 22976
rect 11612 22933 11621 22967
rect 11621 22933 11655 22967
rect 11655 22933 11664 22967
rect 11612 22924 11664 22933
rect 12348 22924 12400 22976
rect 12532 22924 12584 22976
rect 18052 22924 18104 22976
rect 18420 22924 18472 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 4620 22763 4672 22772
rect 4620 22729 4629 22763
rect 4629 22729 4663 22763
rect 4663 22729 4672 22763
rect 4620 22720 4672 22729
rect 8760 22720 8812 22772
rect 12164 22720 12216 22772
rect 14280 22763 14332 22772
rect 14280 22729 14289 22763
rect 14289 22729 14323 22763
rect 14323 22729 14332 22763
rect 14280 22720 14332 22729
rect 19340 22720 19392 22772
rect 19800 22763 19852 22772
rect 19800 22729 19809 22763
rect 19809 22729 19843 22763
rect 19843 22729 19852 22763
rect 19800 22720 19852 22729
rect 23940 22720 23992 22772
rect 24124 22763 24176 22772
rect 24124 22729 24133 22763
rect 24133 22729 24167 22763
rect 24167 22729 24176 22763
rect 24124 22720 24176 22729
rect 13636 22652 13688 22704
rect 17960 22652 18012 22704
rect 22652 22695 22704 22704
rect 22652 22661 22686 22695
rect 22686 22661 22704 22695
rect 22652 22652 22704 22661
rect 4620 22584 4672 22636
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 5632 22516 5684 22568
rect 8576 22584 8628 22636
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 10692 22584 10744 22636
rect 12440 22584 12492 22636
rect 12808 22584 12860 22636
rect 18420 22627 18472 22636
rect 18420 22593 18429 22627
rect 18429 22593 18463 22627
rect 18463 22593 18472 22627
rect 18420 22584 18472 22593
rect 18512 22627 18564 22636
rect 18512 22593 18521 22627
rect 18521 22593 18555 22627
rect 18555 22593 18564 22627
rect 18512 22584 18564 22593
rect 18604 22584 18656 22636
rect 11796 22516 11848 22568
rect 14004 22559 14056 22568
rect 14004 22525 14013 22559
rect 14013 22525 14047 22559
rect 14047 22525 14056 22559
rect 14004 22516 14056 22525
rect 20076 22627 20128 22636
rect 20076 22593 20085 22627
rect 20085 22593 20119 22627
rect 20119 22593 20128 22627
rect 20076 22584 20128 22593
rect 21456 22584 21508 22636
rect 24584 22652 24636 22704
rect 23388 22516 23440 22568
rect 24860 22584 24912 22636
rect 20536 22448 20588 22500
rect 10876 22380 10928 22432
rect 11244 22380 11296 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 10692 22219 10744 22228
rect 10692 22185 10701 22219
rect 10701 22185 10735 22219
rect 10735 22185 10744 22219
rect 10692 22176 10744 22185
rect 12440 22219 12492 22228
rect 12440 22185 12449 22219
rect 12449 22185 12483 22219
rect 12483 22185 12492 22219
rect 12440 22176 12492 22185
rect 14648 22176 14700 22228
rect 18696 22219 18748 22228
rect 18696 22185 18705 22219
rect 18705 22185 18739 22219
rect 18739 22185 18748 22219
rect 18696 22176 18748 22185
rect 9772 22083 9824 22092
rect 9772 22049 9781 22083
rect 9781 22049 9815 22083
rect 9815 22049 9824 22083
rect 9772 22040 9824 22049
rect 1216 21972 1268 22024
rect 10876 22015 10928 22024
rect 10876 21981 10885 22015
rect 10885 21981 10919 22015
rect 10919 21981 10928 22015
rect 10876 21972 10928 21981
rect 11888 21972 11940 22024
rect 4620 21836 4672 21888
rect 12532 22040 12584 22092
rect 22100 22040 22152 22092
rect 12164 21972 12216 22024
rect 14004 21972 14056 22024
rect 13544 21947 13596 21956
rect 13544 21913 13562 21947
rect 13562 21913 13596 21947
rect 13544 21904 13596 21913
rect 13728 21904 13780 21956
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 23388 21972 23440 22024
rect 17224 21947 17276 21956
rect 17224 21913 17233 21947
rect 17233 21913 17267 21947
rect 17267 21913 17276 21947
rect 17224 21904 17276 21913
rect 16856 21879 16908 21888
rect 16856 21845 16865 21879
rect 16865 21845 16899 21879
rect 16899 21845 16908 21879
rect 16856 21836 16908 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 12624 21632 12676 21684
rect 11612 21607 11664 21616
rect 11612 21573 11621 21607
rect 11621 21573 11655 21607
rect 11655 21573 11664 21607
rect 11612 21564 11664 21573
rect 10876 21539 10928 21548
rect 10876 21505 10885 21539
rect 10885 21505 10919 21539
rect 10919 21505 10928 21539
rect 10876 21496 10928 21505
rect 11244 21496 11296 21548
rect 11796 21539 11848 21548
rect 11796 21505 11805 21539
rect 11805 21505 11839 21539
rect 11839 21505 11848 21539
rect 11796 21496 11848 21505
rect 11980 21496 12032 21548
rect 12900 21496 12952 21548
rect 13452 21496 13504 21548
rect 12256 21360 12308 21412
rect 10784 21292 10836 21344
rect 12072 21292 12124 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 11888 21131 11940 21140
rect 11888 21097 11897 21131
rect 11897 21097 11931 21131
rect 11931 21097 11940 21131
rect 11888 21088 11940 21097
rect 13728 21088 13780 21140
rect 9404 20952 9456 21004
rect 12164 20995 12216 21004
rect 12164 20961 12173 20995
rect 12173 20961 12207 20995
rect 12207 20961 12216 20995
rect 12164 20952 12216 20961
rect 10784 20927 10836 20936
rect 10784 20893 10818 20927
rect 10818 20893 10836 20927
rect 10784 20884 10836 20893
rect 15752 20952 15804 21004
rect 12440 20859 12492 20868
rect 12440 20825 12474 20859
rect 12474 20825 12492 20859
rect 12440 20816 12492 20825
rect 15568 20927 15620 20936
rect 15568 20893 15577 20927
rect 15577 20893 15611 20927
rect 15611 20893 15620 20927
rect 15568 20884 15620 20893
rect 16396 20816 16448 20868
rect 15016 20791 15068 20800
rect 15016 20757 15025 20791
rect 15025 20757 15059 20791
rect 15059 20757 15068 20791
rect 15016 20748 15068 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 12440 20544 12492 20553
rect 6460 20451 6512 20460
rect 6460 20417 6469 20451
rect 6469 20417 6503 20451
rect 6503 20417 6512 20451
rect 6460 20408 6512 20417
rect 6552 20408 6604 20460
rect 12532 20476 12584 20528
rect 15016 20476 15068 20528
rect 12256 20451 12308 20460
rect 12256 20417 12265 20451
rect 12265 20417 12299 20451
rect 12299 20417 12308 20451
rect 12256 20408 12308 20417
rect 19892 20476 19944 20528
rect 21824 20476 21876 20528
rect 20260 20408 20312 20460
rect 21180 20408 21232 20460
rect 14004 20340 14056 20392
rect 14556 20383 14608 20392
rect 14556 20349 14565 20383
rect 14565 20349 14599 20383
rect 14599 20349 14608 20383
rect 14556 20340 14608 20349
rect 21088 20383 21140 20392
rect 21088 20349 21097 20383
rect 21097 20349 21131 20383
rect 21131 20349 21140 20383
rect 21088 20340 21140 20349
rect 22928 20408 22980 20460
rect 23388 20408 23440 20460
rect 22008 20272 22060 20324
rect 24492 20340 24544 20392
rect 8116 20204 8168 20256
rect 15200 20204 15252 20256
rect 15568 20204 15620 20256
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 21180 20204 21232 20256
rect 21456 20247 21508 20256
rect 21456 20213 21465 20247
rect 21465 20213 21499 20247
rect 21499 20213 21508 20247
rect 21456 20204 21508 20213
rect 22560 20247 22612 20256
rect 22560 20213 22569 20247
rect 22569 20213 22603 20247
rect 22603 20213 22612 20247
rect 22560 20204 22612 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 5632 20043 5684 20052
rect 5632 20009 5641 20043
rect 5641 20009 5675 20043
rect 5675 20009 5684 20043
rect 5632 20000 5684 20009
rect 6552 20000 6604 20052
rect 18144 20000 18196 20052
rect 15568 19932 15620 19984
rect 8116 19907 8168 19916
rect 8116 19873 8125 19907
rect 8125 19873 8159 19907
rect 8159 19873 8168 19907
rect 8116 19864 8168 19873
rect 14556 19907 14608 19916
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 14556 19864 14608 19873
rect 16028 19864 16080 19916
rect 21088 20000 21140 20052
rect 22008 20000 22060 20052
rect 23664 20000 23716 20052
rect 24308 20000 24360 20052
rect 7840 19796 7892 19848
rect 16396 19839 16448 19848
rect 16396 19805 16405 19839
rect 16405 19805 16439 19839
rect 16439 19805 16448 19839
rect 16396 19796 16448 19805
rect 16488 19839 16540 19848
rect 16488 19805 16497 19839
rect 16497 19805 16531 19839
rect 16531 19805 16540 19839
rect 16488 19796 16540 19805
rect 21548 19932 21600 19984
rect 6736 19728 6788 19780
rect 15016 19728 15068 19780
rect 15752 19728 15804 19780
rect 18144 19839 18196 19848
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 18328 19839 18380 19848
rect 18328 19805 18331 19839
rect 18331 19805 18365 19839
rect 18365 19805 18380 19839
rect 19892 19864 19944 19916
rect 22928 19907 22980 19916
rect 22928 19873 22937 19907
rect 22937 19873 22971 19907
rect 22971 19873 22980 19907
rect 22928 19864 22980 19873
rect 18328 19796 18380 19805
rect 18972 19796 19024 19848
rect 21180 19796 21232 19848
rect 21732 19796 21784 19848
rect 23664 19796 23716 19848
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 16304 19660 16356 19712
rect 17408 19703 17460 19712
rect 17408 19669 17417 19703
rect 17417 19669 17451 19703
rect 17451 19669 17460 19703
rect 17408 19660 17460 19669
rect 19984 19728 20036 19780
rect 18144 19660 18196 19712
rect 18328 19660 18380 19712
rect 19432 19660 19484 19712
rect 21364 19703 21416 19712
rect 21364 19669 21373 19703
rect 21373 19669 21407 19703
rect 21407 19669 21416 19703
rect 21364 19660 21416 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 7840 19499 7892 19508
rect 7840 19465 7849 19499
rect 7849 19465 7883 19499
rect 7883 19465 7892 19499
rect 7840 19456 7892 19465
rect 13452 19499 13504 19508
rect 13452 19465 13461 19499
rect 13461 19465 13495 19499
rect 13495 19465 13504 19499
rect 13452 19456 13504 19465
rect 15016 19499 15068 19508
rect 15016 19465 15025 19499
rect 15025 19465 15059 19499
rect 15059 19465 15068 19499
rect 15016 19456 15068 19465
rect 20904 19456 20956 19508
rect 10876 19388 10928 19440
rect 15752 19431 15804 19440
rect 4620 19252 4672 19304
rect 5908 19320 5960 19372
rect 9404 19320 9456 19372
rect 10600 19363 10652 19372
rect 10600 19329 10609 19363
rect 10609 19329 10643 19363
rect 10643 19329 10652 19363
rect 10600 19320 10652 19329
rect 15752 19397 15761 19431
rect 15761 19397 15795 19431
rect 15795 19397 15804 19431
rect 15752 19388 15804 19397
rect 15568 19320 15620 19372
rect 16396 19388 16448 19440
rect 16028 19363 16080 19372
rect 16028 19329 16037 19363
rect 16037 19329 16071 19363
rect 16071 19329 16080 19363
rect 16028 19320 16080 19329
rect 16488 19320 16540 19372
rect 20260 19320 20312 19372
rect 21824 19456 21876 19508
rect 24308 19499 24360 19508
rect 24308 19465 24317 19499
rect 24317 19465 24351 19499
rect 24351 19465 24360 19499
rect 24308 19456 24360 19465
rect 21548 19388 21600 19440
rect 21456 19320 21508 19372
rect 22008 19320 22060 19372
rect 22928 19320 22980 19372
rect 7104 19295 7156 19304
rect 7104 19261 7113 19295
rect 7113 19261 7147 19295
rect 7147 19261 7156 19295
rect 7104 19252 7156 19261
rect 10048 19295 10100 19304
rect 10048 19261 10057 19295
rect 10057 19261 10091 19295
rect 10091 19261 10100 19295
rect 10048 19252 10100 19261
rect 10508 19252 10560 19304
rect 15660 19252 15712 19304
rect 16212 19252 16264 19304
rect 16304 19252 16356 19304
rect 18144 19295 18196 19304
rect 18144 19261 18153 19295
rect 18153 19261 18187 19295
rect 18187 19261 18196 19295
rect 18144 19252 18196 19261
rect 20352 19295 20404 19304
rect 20352 19261 20361 19295
rect 20361 19261 20395 19295
rect 20395 19261 20404 19295
rect 20352 19252 20404 19261
rect 22376 19295 22428 19304
rect 22376 19261 22385 19295
rect 22385 19261 22419 19295
rect 22419 19261 22428 19295
rect 22376 19252 22428 19261
rect 23848 19295 23900 19304
rect 23848 19261 23857 19295
rect 23857 19261 23891 19295
rect 23891 19261 23900 19295
rect 23848 19252 23900 19261
rect 16672 19184 16724 19236
rect 5448 19159 5500 19168
rect 5448 19125 5457 19159
rect 5457 19125 5491 19159
rect 5491 19125 5500 19159
rect 5448 19116 5500 19125
rect 9220 19116 9272 19168
rect 15844 19159 15896 19168
rect 15844 19125 15853 19159
rect 15853 19125 15887 19159
rect 15887 19125 15896 19159
rect 15844 19116 15896 19125
rect 20996 19116 21048 19168
rect 23112 19116 23164 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 7104 18912 7156 18964
rect 9956 18912 10008 18964
rect 10508 18955 10560 18964
rect 10508 18921 10517 18955
rect 10517 18921 10551 18955
rect 10551 18921 10560 18955
rect 10508 18912 10560 18921
rect 18328 18912 18380 18964
rect 18972 18955 19024 18964
rect 18972 18921 18981 18955
rect 18981 18921 19015 18955
rect 19015 18921 19024 18955
rect 18972 18912 19024 18921
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 20352 18912 20404 18964
rect 21732 18955 21784 18964
rect 21732 18921 21741 18955
rect 21741 18921 21775 18955
rect 21775 18921 21784 18955
rect 21732 18912 21784 18921
rect 21916 18912 21968 18964
rect 23848 18912 23900 18964
rect 9036 18844 9088 18896
rect 9312 18844 9364 18896
rect 10876 18819 10928 18828
rect 10876 18785 10885 18819
rect 10885 18785 10919 18819
rect 10919 18785 10928 18819
rect 10876 18776 10928 18785
rect 24676 18844 24728 18896
rect 15844 18776 15896 18828
rect 20260 18776 20312 18828
rect 24032 18776 24084 18828
rect 24492 18819 24544 18828
rect 24492 18785 24501 18819
rect 24501 18785 24535 18819
rect 24535 18785 24544 18819
rect 24492 18776 24544 18785
rect 3792 18708 3844 18760
rect 4620 18708 4672 18760
rect 5264 18751 5316 18760
rect 5264 18717 5273 18751
rect 5273 18717 5307 18751
rect 5307 18717 5316 18751
rect 5264 18708 5316 18717
rect 7564 18708 7616 18760
rect 9036 18751 9088 18760
rect 9036 18717 9045 18751
rect 9045 18717 9079 18751
rect 9079 18717 9088 18751
rect 9036 18708 9088 18717
rect 9220 18751 9272 18760
rect 9220 18717 9229 18751
rect 9229 18717 9263 18751
rect 9263 18717 9272 18751
rect 9220 18708 9272 18717
rect 5540 18683 5592 18692
rect 5540 18649 5574 18683
rect 5574 18649 5592 18683
rect 5540 18640 5592 18649
rect 6920 18683 6972 18692
rect 6920 18649 6929 18683
rect 6929 18649 6963 18683
rect 6963 18649 6972 18683
rect 6920 18640 6972 18649
rect 4804 18572 4856 18624
rect 6644 18615 6696 18624
rect 6644 18581 6653 18615
rect 6653 18581 6687 18615
rect 6687 18581 6696 18615
rect 6644 18572 6696 18581
rect 6736 18572 6788 18624
rect 7104 18615 7156 18624
rect 7104 18581 7113 18615
rect 7113 18581 7147 18615
rect 7147 18581 7156 18615
rect 7104 18572 7156 18581
rect 7840 18640 7892 18692
rect 9588 18708 9640 18760
rect 9956 18708 10008 18760
rect 18144 18708 18196 18760
rect 18604 18708 18656 18760
rect 17408 18640 17460 18692
rect 9404 18572 9456 18624
rect 10692 18572 10744 18624
rect 10968 18615 11020 18624
rect 10968 18581 10977 18615
rect 10977 18581 11011 18615
rect 11011 18581 11020 18615
rect 10968 18572 11020 18581
rect 17316 18615 17368 18624
rect 17316 18581 17325 18615
rect 17325 18581 17359 18615
rect 17359 18581 17368 18615
rect 17316 18572 17368 18581
rect 20168 18708 20220 18760
rect 23112 18751 23164 18760
rect 23112 18717 23130 18751
rect 23130 18717 23164 18751
rect 23112 18708 23164 18717
rect 23664 18751 23716 18760
rect 23664 18717 23673 18751
rect 23673 18717 23707 18751
rect 23707 18717 23716 18751
rect 23664 18708 23716 18717
rect 20812 18640 20864 18692
rect 24860 18640 24912 18692
rect 20720 18572 20772 18624
rect 21916 18572 21968 18624
rect 23848 18615 23900 18624
rect 23848 18581 23857 18615
rect 23857 18581 23891 18615
rect 23891 18581 23900 18615
rect 23848 18572 23900 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 3792 18411 3844 18420
rect 3792 18377 3801 18411
rect 3801 18377 3835 18411
rect 3835 18377 3844 18411
rect 3792 18368 3844 18377
rect 7104 18368 7156 18420
rect 7840 18411 7892 18420
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 9404 18411 9456 18420
rect 9404 18377 9413 18411
rect 9413 18377 9447 18411
rect 9447 18377 9456 18411
rect 9404 18368 9456 18377
rect 5264 18300 5316 18352
rect 5448 18232 5500 18284
rect 9588 18300 9640 18352
rect 16212 18343 16264 18352
rect 16212 18309 16239 18343
rect 16239 18309 16264 18343
rect 16212 18300 16264 18309
rect 16396 18343 16448 18352
rect 16396 18309 16405 18343
rect 16405 18309 16439 18343
rect 16439 18309 16448 18343
rect 16396 18300 16448 18309
rect 16672 18300 16724 18352
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 7012 18232 7064 18284
rect 11336 18232 11388 18284
rect 8208 18164 8260 18216
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 4712 18096 4764 18148
rect 10048 18096 10100 18148
rect 15384 18164 15436 18216
rect 15660 18232 15712 18284
rect 20812 18411 20864 18420
rect 20812 18377 20821 18411
rect 20821 18377 20855 18411
rect 20855 18377 20864 18411
rect 20812 18368 20864 18377
rect 22376 18411 22428 18420
rect 22376 18377 22385 18411
rect 22385 18377 22419 18411
rect 22419 18377 22428 18411
rect 22376 18368 22428 18377
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 20168 18232 20220 18284
rect 20996 18275 21048 18284
rect 20996 18241 21005 18275
rect 21005 18241 21039 18275
rect 21039 18241 21048 18275
rect 20996 18232 21048 18241
rect 21364 18232 21416 18284
rect 21824 18232 21876 18284
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 22560 18232 22612 18284
rect 23940 18232 23992 18284
rect 24032 18275 24084 18284
rect 24032 18241 24041 18275
rect 24041 18241 24075 18275
rect 24075 18241 24084 18275
rect 24032 18232 24084 18241
rect 16304 18164 16356 18216
rect 16764 18164 16816 18216
rect 21088 18164 21140 18216
rect 16856 18096 16908 18148
rect 18052 18096 18104 18148
rect 848 18028 900 18080
rect 7564 18028 7616 18080
rect 10140 18071 10192 18080
rect 10140 18037 10149 18071
rect 10149 18037 10183 18071
rect 10183 18037 10192 18071
rect 10140 18028 10192 18037
rect 11796 18028 11848 18080
rect 16028 18071 16080 18080
rect 16028 18037 16037 18071
rect 16037 18037 16071 18071
rect 16071 18037 16080 18071
rect 16028 18028 16080 18037
rect 16764 18028 16816 18080
rect 22652 18071 22704 18080
rect 22652 18037 22661 18071
rect 22661 18037 22695 18071
rect 22695 18037 22704 18071
rect 22652 18028 22704 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 7196 17824 7248 17876
rect 8208 17867 8260 17876
rect 8208 17833 8217 17867
rect 8217 17833 8251 17867
rect 8251 17833 8260 17867
rect 8208 17824 8260 17833
rect 9496 17824 9548 17876
rect 10600 17824 10652 17876
rect 11612 17824 11664 17876
rect 16764 17867 16816 17876
rect 16764 17833 16773 17867
rect 16773 17833 16807 17867
rect 16807 17833 16816 17867
rect 16764 17824 16816 17833
rect 20720 17824 20772 17876
rect 23940 17824 23992 17876
rect 24860 17867 24912 17876
rect 24860 17833 24869 17867
rect 24869 17833 24903 17867
rect 24903 17833 24912 17867
rect 24860 17824 24912 17833
rect 4620 17756 4672 17808
rect 12440 17756 12492 17808
rect 20904 17756 20956 17808
rect 9404 17688 9456 17740
rect 17316 17731 17368 17740
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 4804 17552 4856 17604
rect 5264 17620 5316 17672
rect 8024 17620 8076 17672
rect 9312 17663 9364 17672
rect 9312 17629 9321 17663
rect 9321 17629 9355 17663
rect 9355 17629 9364 17663
rect 9312 17620 9364 17629
rect 9496 17663 9548 17672
rect 9496 17629 9505 17663
rect 9505 17629 9539 17663
rect 9539 17629 9548 17663
rect 9496 17620 9548 17629
rect 11796 17620 11848 17672
rect 11888 17663 11940 17672
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 12256 17620 12308 17672
rect 14740 17620 14792 17672
rect 15200 17620 15252 17672
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 15844 17620 15896 17672
rect 17316 17697 17325 17731
rect 17325 17697 17359 17731
rect 17359 17697 17368 17731
rect 17316 17688 17368 17697
rect 3424 17484 3476 17536
rect 4620 17484 4672 17536
rect 6092 17552 6144 17604
rect 17224 17620 17276 17672
rect 20628 17688 20680 17740
rect 17960 17663 18012 17672
rect 17960 17629 17970 17663
rect 17970 17629 18004 17663
rect 18004 17629 18012 17663
rect 17960 17620 18012 17629
rect 18328 17663 18380 17672
rect 18328 17629 18342 17663
rect 18342 17629 18376 17663
rect 18376 17629 18380 17663
rect 18328 17620 18380 17629
rect 5908 17484 5960 17536
rect 9496 17484 9548 17536
rect 18236 17595 18288 17604
rect 18236 17561 18245 17595
rect 18245 17561 18279 17595
rect 18279 17561 18288 17595
rect 18236 17552 18288 17561
rect 22652 17688 22704 17740
rect 23664 17688 23716 17740
rect 23940 17688 23992 17740
rect 21088 17620 21140 17672
rect 21456 17620 21508 17672
rect 20352 17595 20404 17604
rect 20352 17561 20361 17595
rect 20361 17561 20395 17595
rect 20395 17561 20404 17595
rect 20352 17552 20404 17561
rect 21732 17663 21784 17672
rect 21732 17629 21741 17663
rect 21741 17629 21775 17663
rect 21775 17629 21784 17663
rect 21732 17620 21784 17629
rect 21824 17663 21876 17672
rect 21824 17629 21833 17663
rect 21833 17629 21867 17663
rect 21867 17629 21876 17663
rect 21824 17620 21876 17629
rect 21916 17663 21968 17672
rect 21916 17629 21925 17663
rect 21925 17629 21959 17663
rect 21959 17629 21968 17663
rect 21916 17620 21968 17629
rect 22192 17620 22244 17672
rect 24676 17663 24728 17672
rect 24676 17629 24685 17663
rect 24685 17629 24719 17663
rect 24719 17629 24728 17663
rect 24676 17620 24728 17629
rect 20536 17484 20588 17536
rect 23112 17484 23164 17536
rect 23480 17484 23532 17536
rect 23848 17484 23900 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 3148 17280 3200 17332
rect 5540 17280 5592 17332
rect 6092 17323 6144 17332
rect 6092 17289 6101 17323
rect 6101 17289 6135 17323
rect 6135 17289 6144 17323
rect 6092 17280 6144 17289
rect 6920 17280 6972 17332
rect 7288 17280 7340 17332
rect 9588 17280 9640 17332
rect 11704 17280 11756 17332
rect 12164 17280 12216 17332
rect 15844 17323 15896 17332
rect 15844 17289 15853 17323
rect 15853 17289 15887 17323
rect 15887 17289 15896 17323
rect 15844 17280 15896 17289
rect 17960 17280 18012 17332
rect 18052 17323 18104 17332
rect 18052 17289 18061 17323
rect 18061 17289 18095 17323
rect 18095 17289 18104 17323
rect 18052 17280 18104 17289
rect 1308 17144 1360 17196
rect 4620 17212 4672 17264
rect 3424 17144 3476 17196
rect 8024 17212 8076 17264
rect 5632 17076 5684 17128
rect 5908 17187 5960 17196
rect 5908 17153 5917 17187
rect 5917 17153 5951 17187
rect 5951 17153 5960 17187
rect 5908 17144 5960 17153
rect 6644 17144 6696 17196
rect 10140 17212 10192 17264
rect 15384 17212 15436 17264
rect 8208 17144 8260 17196
rect 9404 17144 9456 17196
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 15292 17144 15344 17196
rect 18236 17212 18288 17264
rect 20352 17280 20404 17332
rect 20536 17280 20588 17332
rect 21272 17280 21324 17332
rect 21824 17280 21876 17332
rect 17224 17144 17276 17196
rect 17408 17187 17460 17196
rect 17408 17153 17417 17187
rect 17417 17153 17451 17187
rect 17451 17153 17460 17187
rect 17408 17144 17460 17153
rect 20628 17187 20680 17196
rect 20628 17153 20667 17187
rect 20667 17153 20680 17187
rect 20628 17144 20680 17153
rect 20904 17144 20956 17196
rect 21916 17144 21968 17196
rect 23112 17187 23164 17196
rect 23112 17153 23121 17187
rect 23121 17153 23155 17187
rect 23155 17153 23164 17187
rect 23112 17144 23164 17153
rect 23664 17144 23716 17196
rect 27528 17144 27580 17196
rect 18328 17076 18380 17128
rect 20168 17119 20220 17128
rect 20168 17085 20177 17119
rect 20177 17085 20211 17119
rect 20211 17085 20220 17119
rect 20168 17076 20220 17085
rect 22192 17119 22244 17128
rect 22192 17085 22201 17119
rect 22201 17085 22235 17119
rect 22235 17085 22244 17119
rect 22192 17076 22244 17085
rect 24308 17119 24360 17128
rect 24308 17085 24317 17119
rect 24317 17085 24351 17119
rect 24351 17085 24360 17119
rect 24308 17076 24360 17085
rect 28264 17119 28316 17128
rect 28264 17085 28273 17119
rect 28273 17085 28307 17119
rect 28307 17085 28316 17119
rect 28264 17076 28316 17085
rect 4712 16983 4764 16992
rect 4712 16949 4721 16983
rect 4721 16949 4755 16983
rect 4755 16949 4764 16983
rect 4712 16940 4764 16949
rect 13268 16940 13320 16992
rect 22836 16983 22888 16992
rect 22836 16949 22845 16983
rect 22845 16949 22879 16983
rect 22879 16949 22888 16983
rect 22836 16940 22888 16949
rect 23480 16940 23532 16992
rect 24952 16983 25004 16992
rect 24952 16949 24961 16983
rect 24961 16949 24995 16983
rect 24995 16949 25004 16983
rect 24952 16940 25004 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 4712 16736 4764 16788
rect 8208 16736 8260 16788
rect 24308 16736 24360 16788
rect 10968 16668 11020 16720
rect 7104 16600 7156 16652
rect 5632 16532 5684 16584
rect 7196 16575 7248 16584
rect 7196 16541 7205 16575
rect 7205 16541 7239 16575
rect 7239 16541 7248 16575
rect 7196 16532 7248 16541
rect 7288 16575 7340 16584
rect 7288 16541 7297 16575
rect 7297 16541 7331 16575
rect 7331 16541 7340 16575
rect 7288 16532 7340 16541
rect 7840 16600 7892 16652
rect 11888 16668 11940 16720
rect 11704 16600 11756 16652
rect 12532 16643 12584 16652
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 11888 16532 11940 16584
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 22836 16600 22888 16652
rect 24032 16600 24084 16652
rect 27528 16779 27580 16788
rect 27528 16745 27537 16779
rect 27537 16745 27571 16779
rect 27571 16745 27580 16779
rect 27528 16736 27580 16745
rect 12440 16532 12492 16541
rect 12256 16464 12308 16516
rect 23480 16575 23532 16584
rect 23480 16541 23489 16575
rect 23489 16541 23523 16575
rect 23523 16541 23532 16575
rect 23480 16532 23532 16541
rect 23940 16532 23992 16584
rect 24952 16575 25004 16584
rect 24952 16541 24986 16575
rect 24986 16541 25004 16575
rect 24952 16532 25004 16541
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 13176 16396 13228 16448
rect 23664 16396 23716 16448
rect 27068 16396 27120 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 12532 16192 12584 16244
rect 13636 16192 13688 16244
rect 11796 16099 11848 16108
rect 11796 16065 11805 16099
rect 11805 16065 11839 16099
rect 11839 16065 11848 16099
rect 11796 16056 11848 16065
rect 11888 16031 11940 16040
rect 11888 15997 11897 16031
rect 11897 15997 11931 16031
rect 11931 15997 11940 16031
rect 11888 15988 11940 15997
rect 13176 16099 13228 16108
rect 13176 16065 13185 16099
rect 13185 16065 13219 16099
rect 13219 16065 13228 16099
rect 13176 16056 13228 16065
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 13912 16099 13964 16108
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 15292 16124 15344 16176
rect 14280 16056 14332 16108
rect 27068 16099 27120 16108
rect 27068 16065 27077 16099
rect 27077 16065 27111 16099
rect 27111 16065 27120 16099
rect 27068 16056 27120 16065
rect 28264 16031 28316 16040
rect 28264 15997 28273 16031
rect 28273 15997 28307 16031
rect 28307 15997 28316 16031
rect 28264 15988 28316 15997
rect 15752 15920 15804 15972
rect 14464 15852 14516 15904
rect 14740 15895 14792 15904
rect 14740 15861 14749 15895
rect 14749 15861 14783 15895
rect 14783 15861 14792 15895
rect 14740 15852 14792 15861
rect 23940 15852 23992 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 12440 15648 12492 15700
rect 13636 15691 13688 15700
rect 13636 15657 13645 15691
rect 13645 15657 13679 15691
rect 13679 15657 13688 15691
rect 13636 15648 13688 15657
rect 14832 15691 14884 15700
rect 14832 15657 14841 15691
rect 14841 15657 14875 15691
rect 14875 15657 14884 15691
rect 14832 15648 14884 15657
rect 12256 15512 12308 15564
rect 9772 15444 9824 15496
rect 11704 15444 11756 15496
rect 12716 15487 12768 15496
rect 12716 15453 12725 15487
rect 12725 15453 12759 15487
rect 12759 15453 12768 15487
rect 12716 15444 12768 15453
rect 14740 15512 14792 15564
rect 13636 15444 13688 15496
rect 10968 15419 11020 15428
rect 10968 15385 11002 15419
rect 11002 15385 11020 15419
rect 10968 15376 11020 15385
rect 13820 15376 13872 15428
rect 13912 15308 13964 15360
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 15660 15419 15712 15428
rect 15660 15385 15669 15419
rect 15669 15385 15703 15419
rect 15703 15385 15712 15419
rect 15660 15376 15712 15385
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 10968 15104 11020 15156
rect 13820 15104 13872 15156
rect 15292 15104 15344 15156
rect 9772 14968 9824 15020
rect 11612 14968 11664 15020
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 14832 14968 14884 15020
rect 16580 14968 16632 15020
rect 25136 14968 25188 15020
rect 9680 14900 9732 14952
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 14464 14943 14516 14952
rect 14464 14909 14473 14943
rect 14473 14909 14507 14943
rect 14507 14909 14516 14943
rect 14464 14900 14516 14909
rect 14924 14943 14976 14952
rect 14924 14909 14933 14943
rect 14933 14909 14967 14943
rect 14967 14909 14976 14943
rect 14924 14900 14976 14909
rect 25412 14900 25464 14952
rect 12992 14807 13044 14816
rect 12992 14773 13001 14807
rect 13001 14773 13035 14807
rect 13035 14773 13044 14807
rect 12992 14764 13044 14773
rect 15568 14764 15620 14816
rect 23664 14807 23716 14816
rect 23664 14773 23673 14807
rect 23673 14773 23707 14807
rect 23707 14773 23716 14807
rect 23664 14764 23716 14773
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 8484 14603 8536 14612
rect 8484 14569 8493 14603
rect 8493 14569 8527 14603
rect 8527 14569 8536 14603
rect 8484 14560 8536 14569
rect 9772 14603 9824 14612
rect 9772 14569 9781 14603
rect 9781 14569 9815 14603
rect 9815 14569 9824 14603
rect 9772 14560 9824 14569
rect 11336 14603 11388 14612
rect 11336 14569 11345 14603
rect 11345 14569 11379 14603
rect 11379 14569 11388 14603
rect 11336 14560 11388 14569
rect 11888 14560 11940 14612
rect 14372 14560 14424 14612
rect 14924 14560 14976 14612
rect 25136 14603 25188 14612
rect 25136 14569 25145 14603
rect 25145 14569 25179 14603
rect 25179 14569 25188 14603
rect 25136 14560 25188 14569
rect 25412 14603 25464 14612
rect 25412 14569 25421 14603
rect 25421 14569 25455 14603
rect 25455 14569 25464 14603
rect 25412 14560 25464 14569
rect 12532 14492 12584 14544
rect 7104 14424 7156 14476
rect 7380 14288 7432 14340
rect 7932 14399 7984 14408
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 12716 14424 12768 14476
rect 11336 14356 11388 14408
rect 14280 14356 14332 14408
rect 14372 14356 14424 14408
rect 15384 14399 15436 14408
rect 15384 14365 15393 14399
rect 15393 14365 15427 14399
rect 15427 14365 15436 14399
rect 15384 14356 15436 14365
rect 15568 14399 15620 14408
rect 15568 14365 15577 14399
rect 15577 14365 15611 14399
rect 15611 14365 15620 14399
rect 15568 14356 15620 14365
rect 19616 14356 19668 14408
rect 20168 14356 20220 14408
rect 7564 14263 7616 14272
rect 7564 14229 7573 14263
rect 7573 14229 7607 14263
rect 7607 14229 7616 14263
rect 7564 14220 7616 14229
rect 8300 14288 8352 14340
rect 20260 14288 20312 14340
rect 9680 14220 9732 14272
rect 20628 14220 20680 14272
rect 24124 14356 24176 14408
rect 24860 14356 24912 14408
rect 28448 14399 28500 14408
rect 28448 14365 28457 14399
rect 28457 14365 28491 14399
rect 28491 14365 28500 14399
rect 28448 14356 28500 14365
rect 23204 14288 23256 14340
rect 21640 14263 21692 14272
rect 21640 14229 21649 14263
rect 21649 14229 21683 14263
rect 21683 14229 21692 14263
rect 21640 14220 21692 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 7932 14016 7984 14068
rect 14372 14059 14424 14068
rect 14372 14025 14381 14059
rect 14381 14025 14415 14059
rect 14415 14025 14424 14059
rect 14372 14016 14424 14025
rect 15292 14016 15344 14068
rect 20260 14059 20312 14068
rect 20260 14025 20269 14059
rect 20269 14025 20303 14059
rect 20303 14025 20312 14059
rect 20260 14016 20312 14025
rect 23204 14059 23256 14068
rect 23204 14025 23213 14059
rect 23213 14025 23247 14059
rect 23247 14025 23256 14059
rect 23204 14016 23256 14025
rect 7104 13812 7156 13864
rect 8116 13855 8168 13864
rect 8116 13821 8125 13855
rect 8125 13821 8159 13855
rect 8159 13821 8168 13855
rect 8116 13812 8168 13821
rect 10140 13923 10192 13932
rect 10140 13889 10149 13923
rect 10149 13889 10183 13923
rect 10183 13889 10192 13923
rect 10140 13880 10192 13889
rect 10324 13812 10376 13864
rect 10600 13880 10652 13932
rect 12440 13880 12492 13932
rect 13544 13880 13596 13932
rect 14924 13880 14976 13932
rect 20444 13948 20496 14000
rect 10968 13812 11020 13864
rect 12900 13744 12952 13796
rect 17408 13744 17460 13796
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 20536 13880 20588 13889
rect 20812 13923 20864 13932
rect 20812 13889 20821 13923
rect 20821 13889 20855 13923
rect 20855 13889 20864 13923
rect 20812 13880 20864 13889
rect 24952 13880 25004 13932
rect 19984 13744 20036 13796
rect 23756 13855 23808 13864
rect 23756 13821 23765 13855
rect 23765 13821 23799 13855
rect 23799 13821 23808 13855
rect 23756 13812 23808 13821
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 10232 13676 10284 13728
rect 24216 13719 24268 13728
rect 24216 13685 24225 13719
rect 24225 13685 24259 13719
rect 24259 13685 24268 13719
rect 24216 13676 24268 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 8116 13515 8168 13524
rect 8116 13481 8125 13515
rect 8125 13481 8159 13515
rect 8159 13481 8168 13515
rect 8116 13472 8168 13481
rect 9772 13472 9824 13524
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 10324 13515 10376 13524
rect 10324 13481 10333 13515
rect 10333 13481 10367 13515
rect 10367 13481 10376 13515
rect 10324 13472 10376 13481
rect 12716 13472 12768 13524
rect 13544 13515 13596 13524
rect 13544 13481 13553 13515
rect 13553 13481 13587 13515
rect 13587 13481 13596 13515
rect 13544 13472 13596 13481
rect 15660 13404 15712 13456
rect 10600 13379 10652 13388
rect 10600 13345 10609 13379
rect 10609 13345 10643 13379
rect 10643 13345 10652 13379
rect 10600 13336 10652 13345
rect 16580 13379 16632 13388
rect 16580 13345 16589 13379
rect 16589 13345 16623 13379
rect 16623 13345 16632 13379
rect 16580 13336 16632 13345
rect 7288 13268 7340 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9588 13268 9640 13320
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 11336 13268 11388 13320
rect 12992 13268 13044 13320
rect 17224 13336 17276 13388
rect 24400 13404 24452 13456
rect 21732 13336 21784 13388
rect 7012 13243 7064 13252
rect 7012 13209 7046 13243
rect 7046 13209 7064 13243
rect 7012 13200 7064 13209
rect 10876 13243 10928 13252
rect 10876 13209 10910 13243
rect 10910 13209 10928 13243
rect 10876 13200 10928 13209
rect 9956 13175 10008 13184
rect 9956 13141 9965 13175
rect 9965 13141 9999 13175
rect 9999 13141 10008 13175
rect 9956 13132 10008 13141
rect 10140 13132 10192 13184
rect 16856 13268 16908 13320
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 19432 13268 19484 13320
rect 20076 13311 20128 13320
rect 20076 13277 20085 13311
rect 20085 13277 20119 13311
rect 20119 13277 20128 13311
rect 20076 13268 20128 13277
rect 15200 13132 15252 13184
rect 16304 13175 16356 13184
rect 16304 13141 16313 13175
rect 16313 13141 16347 13175
rect 16347 13141 16356 13175
rect 16304 13132 16356 13141
rect 19340 13132 19392 13184
rect 19708 13175 19760 13184
rect 19708 13141 19717 13175
rect 19717 13141 19751 13175
rect 19751 13141 19760 13175
rect 19708 13132 19760 13141
rect 19984 13243 20036 13252
rect 19984 13209 19993 13243
rect 19993 13209 20027 13243
rect 20027 13209 20036 13243
rect 19984 13200 20036 13209
rect 20628 13311 20680 13320
rect 20628 13277 20636 13311
rect 20636 13277 20670 13311
rect 20670 13277 20680 13311
rect 20628 13268 20680 13277
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 23664 13268 23716 13320
rect 23020 13132 23072 13184
rect 23664 13132 23716 13184
rect 23940 13132 23992 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 8392 12928 8444 12980
rect 5540 12792 5592 12844
rect 6920 12860 6972 12912
rect 6092 12767 6144 12776
rect 6092 12733 6101 12767
rect 6101 12733 6135 12767
rect 6135 12733 6144 12767
rect 6092 12724 6144 12733
rect 7380 12860 7432 12912
rect 7564 12903 7616 12912
rect 7564 12869 7598 12903
rect 7598 12869 7616 12903
rect 7564 12860 7616 12869
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 9128 12928 9180 12980
rect 10876 12971 10928 12980
rect 10876 12937 10885 12971
rect 10885 12937 10919 12971
rect 10919 12937 10928 12971
rect 10876 12928 10928 12937
rect 11336 12928 11388 12980
rect 9956 12860 10008 12912
rect 12900 12928 12952 12980
rect 20536 12928 20588 12980
rect 20628 12928 20680 12980
rect 23572 12928 23624 12980
rect 24860 12928 24912 12980
rect 24952 12971 25004 12980
rect 24952 12937 24961 12971
rect 24961 12937 24995 12971
rect 24995 12937 25004 12971
rect 24952 12928 25004 12937
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 11612 12767 11664 12776
rect 11612 12733 11621 12767
rect 11621 12733 11655 12767
rect 11655 12733 11664 12767
rect 11612 12724 11664 12733
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 15660 12792 15712 12844
rect 19984 12860 20036 12912
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 12624 12767 12676 12776
rect 12624 12733 12633 12767
rect 12633 12733 12667 12767
rect 12667 12733 12676 12767
rect 12624 12724 12676 12733
rect 16304 12724 16356 12776
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 18512 12835 18564 12844
rect 18512 12801 18521 12835
rect 18521 12801 18555 12835
rect 18555 12801 18564 12835
rect 18512 12792 18564 12801
rect 23756 12903 23808 12912
rect 23756 12869 23765 12903
rect 23765 12869 23799 12903
rect 23799 12869 23808 12903
rect 23756 12860 23808 12869
rect 24216 12903 24268 12912
rect 24216 12869 24225 12903
rect 24225 12869 24259 12903
rect 24259 12869 24268 12903
rect 24216 12860 24268 12869
rect 17408 12767 17460 12776
rect 17408 12733 17417 12767
rect 17417 12733 17451 12767
rect 17451 12733 17460 12767
rect 17408 12724 17460 12733
rect 19340 12767 19392 12776
rect 19340 12733 19349 12767
rect 19349 12733 19383 12767
rect 19383 12733 19392 12767
rect 19340 12724 19392 12733
rect 21272 12835 21324 12844
rect 21272 12801 21281 12835
rect 21281 12801 21315 12835
rect 21315 12801 21324 12835
rect 21272 12792 21324 12801
rect 21640 12792 21692 12844
rect 20076 12767 20128 12776
rect 20076 12733 20085 12767
rect 20085 12733 20119 12767
rect 20119 12733 20128 12767
rect 20076 12724 20128 12733
rect 16672 12656 16724 12708
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 17224 12656 17276 12708
rect 19432 12656 19484 12708
rect 21732 12724 21784 12776
rect 21824 12724 21876 12776
rect 20904 12699 20956 12708
rect 20904 12665 20913 12699
rect 20913 12665 20947 12699
rect 20947 12665 20956 12699
rect 20904 12656 20956 12665
rect 22468 12792 22520 12844
rect 23664 12792 23716 12844
rect 24032 12792 24084 12844
rect 23020 12767 23072 12776
rect 23020 12733 23029 12767
rect 23029 12733 23063 12767
rect 23063 12733 23072 12767
rect 23020 12724 23072 12733
rect 23480 12699 23532 12708
rect 23480 12665 23489 12699
rect 23489 12665 23523 12699
rect 23523 12665 23532 12699
rect 23480 12656 23532 12665
rect 24584 12835 24636 12844
rect 24584 12801 24593 12835
rect 24593 12801 24627 12835
rect 24627 12801 24636 12835
rect 24584 12792 24636 12801
rect 24768 12835 24820 12844
rect 24768 12801 24777 12835
rect 24777 12801 24811 12835
rect 24811 12801 24820 12835
rect 24768 12792 24820 12801
rect 17408 12588 17460 12640
rect 18236 12631 18288 12640
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 9404 12384 9456 12436
rect 11336 12427 11388 12436
rect 11336 12393 11345 12427
rect 11345 12393 11379 12427
rect 11379 12393 11388 12427
rect 11336 12384 11388 12393
rect 11612 12427 11664 12436
rect 11612 12393 11621 12427
rect 11621 12393 11655 12427
rect 11655 12393 11664 12427
rect 11612 12384 11664 12393
rect 12624 12384 12676 12436
rect 14464 12384 14516 12436
rect 16672 12384 16724 12436
rect 16856 12384 16908 12436
rect 18512 12384 18564 12436
rect 18052 12316 18104 12368
rect 16764 12248 16816 12300
rect 5448 12180 5500 12232
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 5724 12112 5776 12164
rect 7932 12112 7984 12164
rect 9956 12223 10008 12232
rect 9956 12189 9965 12223
rect 9965 12189 9999 12223
rect 9999 12189 10008 12223
rect 9956 12180 10008 12189
rect 10600 12180 10652 12232
rect 12440 12180 12492 12232
rect 18236 12248 18288 12300
rect 17960 12180 18012 12232
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 20444 12248 20496 12300
rect 23572 12316 23624 12368
rect 23480 12248 23532 12300
rect 10232 12155 10284 12164
rect 10232 12121 10266 12155
rect 10266 12121 10284 12155
rect 10232 12112 10284 12121
rect 10692 12112 10744 12164
rect 17868 12112 17920 12164
rect 19432 12180 19484 12232
rect 20904 12180 20956 12232
rect 21824 12223 21876 12232
rect 21824 12189 21833 12223
rect 21833 12189 21867 12223
rect 21867 12189 21876 12223
rect 21824 12180 21876 12189
rect 22744 12223 22796 12232
rect 22744 12189 22753 12223
rect 22753 12189 22787 12223
rect 22787 12189 22796 12223
rect 22744 12180 22796 12189
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 10048 12044 10100 12096
rect 16028 12087 16080 12096
rect 16028 12053 16037 12087
rect 16037 12053 16071 12087
rect 16071 12053 16080 12087
rect 16028 12044 16080 12053
rect 16304 12087 16356 12096
rect 16304 12053 16313 12087
rect 16313 12053 16347 12087
rect 16347 12053 16356 12087
rect 16304 12044 16356 12053
rect 22284 12112 22336 12164
rect 20260 12087 20312 12096
rect 20260 12053 20269 12087
rect 20269 12053 20303 12087
rect 20303 12053 20312 12087
rect 20260 12044 20312 12053
rect 21180 12044 21232 12096
rect 21456 12044 21508 12096
rect 22192 12087 22244 12096
rect 22192 12053 22201 12087
rect 22201 12053 22235 12087
rect 22235 12053 22244 12087
rect 22192 12044 22244 12053
rect 25136 12087 25188 12096
rect 25136 12053 25145 12087
rect 25145 12053 25179 12087
rect 25179 12053 25188 12087
rect 25136 12044 25188 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 6092 11840 6144 11892
rect 8300 11840 8352 11892
rect 16856 11840 16908 11892
rect 17592 11883 17644 11892
rect 17592 11849 17601 11883
rect 17601 11849 17635 11883
rect 17635 11849 17644 11883
rect 17592 11840 17644 11849
rect 21824 11840 21876 11892
rect 22468 11883 22520 11892
rect 22468 11849 22477 11883
rect 22477 11849 22511 11883
rect 22511 11849 22520 11883
rect 22468 11840 22520 11849
rect 22744 11883 22796 11892
rect 22744 11849 22753 11883
rect 22753 11849 22787 11883
rect 22787 11849 22796 11883
rect 22744 11840 22796 11849
rect 5540 11747 5592 11756
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 5908 11704 5960 11756
rect 8300 11747 8352 11756
rect 8300 11713 8309 11747
rect 8309 11713 8343 11747
rect 8343 11713 8352 11747
rect 8300 11704 8352 11713
rect 9864 11704 9916 11756
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 11336 11704 11388 11756
rect 14372 11747 14424 11756
rect 14372 11713 14381 11747
rect 14381 11713 14415 11747
rect 14415 11713 14424 11747
rect 14372 11704 14424 11713
rect 14464 11704 14516 11756
rect 15200 11704 15252 11756
rect 6828 11636 6880 11688
rect 8484 11636 8536 11688
rect 14280 11636 14332 11688
rect 14924 11636 14976 11688
rect 16304 11704 16356 11756
rect 18144 11772 18196 11824
rect 21272 11772 21324 11824
rect 24768 11840 24820 11892
rect 16580 11636 16632 11688
rect 17868 11704 17920 11756
rect 19892 11747 19944 11756
rect 19892 11713 19926 11747
rect 19926 11713 19944 11747
rect 19892 11704 19944 11713
rect 21456 11747 21508 11756
rect 21456 11713 21465 11747
rect 21465 11713 21499 11747
rect 21499 11713 21508 11747
rect 21456 11704 21508 11713
rect 21732 11704 21784 11756
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 19616 11679 19668 11688
rect 19616 11645 19625 11679
rect 19625 11645 19659 11679
rect 19659 11645 19668 11679
rect 19616 11636 19668 11645
rect 24124 11747 24176 11756
rect 24124 11713 24133 11747
rect 24133 11713 24167 11747
rect 24167 11713 24176 11747
rect 24124 11704 24176 11713
rect 25136 11747 25188 11756
rect 25136 11713 25145 11747
rect 25145 11713 25179 11747
rect 25179 11713 25188 11747
rect 25136 11704 25188 11713
rect 24492 11679 24544 11688
rect 24492 11645 24501 11679
rect 24501 11645 24535 11679
rect 24535 11645 24544 11679
rect 24492 11636 24544 11645
rect 24768 11636 24820 11688
rect 19524 11568 19576 11620
rect 5724 11500 5776 11552
rect 8300 11500 8352 11552
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 14096 11500 14148 11552
rect 15844 11543 15896 11552
rect 15844 11509 15853 11543
rect 15853 11509 15887 11543
rect 15887 11509 15896 11543
rect 15844 11500 15896 11509
rect 17960 11543 18012 11552
rect 17960 11509 17969 11543
rect 17969 11509 18003 11543
rect 18003 11509 18012 11543
rect 17960 11500 18012 11509
rect 20812 11500 20864 11552
rect 22100 11500 22152 11552
rect 24584 11500 24636 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 7932 11339 7984 11348
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 9680 11296 9732 11348
rect 10692 11296 10744 11348
rect 14924 11339 14976 11348
rect 14924 11305 14933 11339
rect 14933 11305 14967 11339
rect 14967 11305 14976 11339
rect 14924 11296 14976 11305
rect 16028 11296 16080 11348
rect 7012 11228 7064 11280
rect 5448 11203 5500 11212
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 8300 11203 8352 11212
rect 8300 11169 8309 11203
rect 8309 11169 8343 11203
rect 8343 11169 8352 11203
rect 8300 11160 8352 11169
rect 10048 11160 10100 11212
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 17960 11296 18012 11348
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 19892 11339 19944 11348
rect 19892 11305 19901 11339
rect 19901 11305 19935 11339
rect 19935 11305 19944 11339
rect 19892 11296 19944 11305
rect 22100 11339 22152 11348
rect 22100 11305 22109 11339
rect 22109 11305 22143 11339
rect 22143 11305 22152 11339
rect 22100 11296 22152 11305
rect 22284 11296 22336 11348
rect 23848 11339 23900 11348
rect 23848 11305 23857 11339
rect 23857 11305 23891 11339
rect 23891 11305 23900 11339
rect 23848 11296 23900 11305
rect 17408 11228 17460 11280
rect 20812 11228 20864 11280
rect 23664 11228 23716 11280
rect 24768 11228 24820 11280
rect 5724 11135 5776 11144
rect 5724 11101 5758 11135
rect 5758 11101 5776 11135
rect 5724 11092 5776 11101
rect 7380 11092 7432 11144
rect 8392 11092 8444 11144
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 9588 11092 9640 11144
rect 16212 11092 16264 11144
rect 19616 11160 19668 11212
rect 20260 11160 20312 11212
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 19524 11092 19576 11144
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 22192 11092 22244 11144
rect 24492 11092 24544 11144
rect 8484 11024 8536 11076
rect 13452 11024 13504 11076
rect 15844 11024 15896 11076
rect 18144 11024 18196 11076
rect 23848 11024 23900 11076
rect 28264 11024 28316 11076
rect 17040 10999 17092 11008
rect 17040 10965 17049 10999
rect 17049 10965 17083 10999
rect 17083 10965 17092 10999
rect 17040 10956 17092 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 9864 10752 9916 10804
rect 13452 10795 13504 10804
rect 13452 10761 13461 10795
rect 13461 10761 13495 10795
rect 13495 10761 13504 10795
rect 13452 10752 13504 10761
rect 14924 10752 14976 10804
rect 18236 10752 18288 10804
rect 19524 10752 19576 10804
rect 15200 10684 15252 10736
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 10600 10616 10652 10668
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 14464 10616 14516 10668
rect 17040 10616 17092 10668
rect 18052 10616 18104 10668
rect 14372 10523 14424 10532
rect 14372 10489 14381 10523
rect 14381 10489 14415 10523
rect 14415 10489 14424 10523
rect 14372 10480 14424 10489
rect 15936 10412 15988 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 18052 10208 18104 10260
rect 16212 10115 16264 10124
rect 16212 10081 16221 10115
rect 16221 10081 16255 10115
rect 16255 10081 16264 10115
rect 16212 10072 16264 10081
rect 15200 10004 15252 10056
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 15752 9664 15804 9716
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 28264 8619 28316 8628
rect 28264 8585 28273 8619
rect 28273 8585 28307 8619
rect 28307 8585 28316 8619
rect 28264 8576 28316 8585
rect 28448 8483 28500 8492
rect 28448 8449 28457 8483
rect 28457 8449 28491 8483
rect 28491 8449 28500 8483
rect 28448 8440 28500 8449
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 28264 8032 28316 8084
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 5908 2635 5960 2644
rect 5908 2601 5917 2635
rect 5917 2601 5951 2635
rect 5951 2601 5960 2635
rect 5908 2592 5960 2601
rect 5816 2388 5868 2440
rect 21916 2388 21968 2440
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5170 49314 5226 50000
rect 21914 49314 21970 50000
rect 24490 49314 24546 50000
rect 5170 49286 5488 49314
rect 5170 49200 5226 49286
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4712 47184 4764 47190
rect 4712 47126 4764 47132
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 110 44568 166 44577
rect 110 44503 166 44512
rect 124 27946 152 44503
rect 4724 44402 4752 47126
rect 5460 47054 5488 49286
rect 21914 49286 22048 49314
rect 21914 49200 21970 49286
rect 22020 47122 22048 49286
rect 24490 49286 24624 49314
rect 24490 49200 24546 49286
rect 24596 47258 24624 49286
rect 24584 47252 24636 47258
rect 24584 47194 24636 47200
rect 22008 47116 22060 47122
rect 22008 47058 22060 47064
rect 5448 47048 5500 47054
rect 5448 46990 5500 46996
rect 22100 47048 22152 47054
rect 22100 46990 22152 46996
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 10048 45552 10100 45558
rect 10048 45494 10100 45500
rect 20628 45552 20680 45558
rect 20628 45494 20680 45500
rect 9956 45348 10008 45354
rect 9956 45290 10008 45296
rect 9404 45280 9456 45286
rect 9404 45222 9456 45228
rect 7472 44872 7524 44878
rect 7472 44814 7524 44820
rect 6920 44736 6972 44742
rect 6920 44678 6972 44684
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 4712 44396 4764 44402
rect 4712 44338 4764 44344
rect 5632 44396 5684 44402
rect 5632 44338 5684 44344
rect 4712 44192 4764 44198
rect 4712 44134 4764 44140
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4528 43784 4580 43790
rect 4580 43732 4660 43738
rect 4528 43726 4660 43732
rect 4540 43710 4660 43726
rect 4724 43722 4752 44134
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4632 42684 4660 43710
rect 4712 43716 4764 43722
rect 4712 43658 4764 43664
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 4712 42696 4764 42702
rect 4632 42656 4712 42684
rect 4712 42638 4764 42644
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4724 41138 4752 42638
rect 5448 42628 5500 42634
rect 5448 42570 5500 42576
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 5460 42362 5488 42570
rect 5448 42356 5500 42362
rect 5448 42298 5500 42304
rect 5644 42226 5672 44338
rect 6932 44198 6960 44678
rect 7196 44328 7248 44334
rect 7196 44270 7248 44276
rect 6920 44192 6972 44198
rect 6920 44134 6972 44140
rect 7208 43790 7236 44270
rect 7484 43994 7512 44814
rect 7840 44736 7892 44742
rect 7840 44678 7892 44684
rect 9220 44736 9272 44742
rect 9220 44678 9272 44684
rect 7472 43988 7524 43994
rect 7472 43930 7524 43936
rect 7196 43784 7248 43790
rect 7196 43726 7248 43732
rect 7852 43722 7880 44678
rect 7932 44192 7984 44198
rect 7932 44134 7984 44140
rect 8576 44192 8628 44198
rect 8576 44134 8628 44140
rect 7840 43716 7892 43722
rect 7840 43658 7892 43664
rect 6460 43648 6512 43654
rect 6460 43590 6512 43596
rect 6472 43314 6500 43590
rect 6460 43308 6512 43314
rect 6460 43250 6512 43256
rect 5816 43104 5868 43110
rect 5816 43046 5868 43052
rect 6828 43104 6880 43110
rect 6828 43046 6880 43052
rect 5828 42226 5856 43046
rect 6460 42560 6512 42566
rect 6460 42502 6512 42508
rect 6472 42226 6500 42502
rect 5632 42220 5684 42226
rect 5632 42162 5684 42168
rect 5816 42220 5868 42226
rect 5816 42162 5868 42168
rect 6460 42220 6512 42226
rect 6460 42162 6512 42168
rect 5644 41614 5672 42162
rect 5632 41608 5684 41614
rect 5632 41550 5684 41556
rect 5540 41472 5592 41478
rect 5540 41414 5592 41420
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 5448 41200 5500 41206
rect 5448 41142 5500 41148
rect 4712 41132 4764 41138
rect 4712 41074 4764 41080
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 5460 39522 5488 41142
rect 5552 41138 5580 41414
rect 5540 41132 5592 41138
rect 5540 41074 5592 41080
rect 5644 40526 5672 41550
rect 6840 41274 6868 43046
rect 7104 42016 7156 42022
rect 7104 41958 7156 41964
rect 7116 41682 7144 41958
rect 7104 41676 7156 41682
rect 7104 41618 7156 41624
rect 6828 41268 6880 41274
rect 6828 41210 6880 41216
rect 6644 41200 6696 41206
rect 6644 41142 6696 41148
rect 6656 40526 6684 41142
rect 6840 40730 6868 41210
rect 7116 41188 7144 41618
rect 7196 41200 7248 41206
rect 7116 41160 7196 41188
rect 6828 40724 6880 40730
rect 6828 40666 6880 40672
rect 7116 40526 7144 41160
rect 7196 41142 7248 41148
rect 7944 41138 7972 44134
rect 7932 41132 7984 41138
rect 7932 41074 7984 41080
rect 7472 40928 7524 40934
rect 7472 40870 7524 40876
rect 5632 40520 5684 40526
rect 5632 40462 5684 40468
rect 6644 40520 6696 40526
rect 6644 40462 6696 40468
rect 7104 40520 7156 40526
rect 7104 40462 7156 40468
rect 7288 40452 7340 40458
rect 7288 40394 7340 40400
rect 5908 40384 5960 40390
rect 5908 40326 5960 40332
rect 5460 39506 5580 39522
rect 5460 39500 5592 39506
rect 5460 39494 5540 39500
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 1216 38344 1268 38350
rect 1216 38286 1268 38292
rect 1228 38185 1256 38286
rect 1676 38208 1728 38214
rect 1214 38176 1270 38185
rect 1676 38150 1728 38156
rect 1214 38111 1270 38120
rect 1688 37874 1716 38150
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 5460 37942 5488 39494
rect 5540 39442 5592 39448
rect 5920 39438 5948 40326
rect 7012 39976 7064 39982
rect 7012 39918 7064 39924
rect 7024 39642 7052 39918
rect 7012 39636 7064 39642
rect 7012 39578 7064 39584
rect 5908 39432 5960 39438
rect 5908 39374 5960 39380
rect 7300 39370 7328 40394
rect 7288 39364 7340 39370
rect 7288 39306 7340 39312
rect 7300 38350 7328 39306
rect 7484 38962 7512 40870
rect 7748 40724 7800 40730
rect 7748 40666 7800 40672
rect 7656 40588 7708 40594
rect 7656 40530 7708 40536
rect 7668 40186 7696 40530
rect 7656 40180 7708 40186
rect 7656 40122 7708 40128
rect 7668 39506 7696 40122
rect 7656 39500 7708 39506
rect 7656 39442 7708 39448
rect 7760 39098 7788 40666
rect 7944 40594 7972 41074
rect 8588 40730 8616 44134
rect 8576 40724 8628 40730
rect 8576 40666 8628 40672
rect 7840 40588 7892 40594
rect 7840 40530 7892 40536
rect 7932 40588 7984 40594
rect 7932 40530 7984 40536
rect 7852 40186 7880 40530
rect 7840 40180 7892 40186
rect 7840 40122 7892 40128
rect 7852 39370 7880 40122
rect 8024 40044 8076 40050
rect 8024 39986 8076 39992
rect 8208 40044 8260 40050
rect 8208 39986 8260 39992
rect 7840 39364 7892 39370
rect 7840 39306 7892 39312
rect 7748 39092 7800 39098
rect 7748 39034 7800 39040
rect 7852 38962 7880 39306
rect 8036 38962 8064 39986
rect 8220 39642 8248 39986
rect 8208 39636 8260 39642
rect 8208 39578 8260 39584
rect 8220 39030 8248 39578
rect 9232 39438 9260 44678
rect 9416 44402 9444 45222
rect 9496 44872 9548 44878
rect 9496 44814 9548 44820
rect 9404 44396 9456 44402
rect 9404 44338 9456 44344
rect 9508 40730 9536 44814
rect 9968 44810 9996 45290
rect 10060 45082 10088 45494
rect 10876 45484 10928 45490
rect 10876 45426 10928 45432
rect 11796 45484 11848 45490
rect 11796 45426 11848 45432
rect 11888 45484 11940 45490
rect 11888 45426 11940 45432
rect 13912 45484 13964 45490
rect 13912 45426 13964 45432
rect 14740 45484 14792 45490
rect 14740 45426 14792 45432
rect 16028 45484 16080 45490
rect 16028 45426 16080 45432
rect 19524 45484 19576 45490
rect 19524 45426 19576 45432
rect 19984 45484 20036 45490
rect 19984 45426 20036 45432
rect 10888 45354 10916 45426
rect 11704 45416 11756 45422
rect 11704 45358 11756 45364
rect 10876 45348 10928 45354
rect 10876 45290 10928 45296
rect 11060 45280 11112 45286
rect 11060 45222 11112 45228
rect 10048 45076 10100 45082
rect 10048 45018 10100 45024
rect 9956 44804 10008 44810
rect 9956 44746 10008 44752
rect 9864 44328 9916 44334
rect 9864 44270 9916 44276
rect 9876 43858 9904 44270
rect 9864 43852 9916 43858
rect 9864 43794 9916 43800
rect 9968 43722 9996 44746
rect 9956 43716 10008 43722
rect 9956 43658 10008 43664
rect 9968 42838 9996 43658
rect 10060 43314 10088 45018
rect 10784 44872 10836 44878
rect 10784 44814 10836 44820
rect 10796 44538 10824 44814
rect 10784 44532 10836 44538
rect 10784 44474 10836 44480
rect 10968 43784 11020 43790
rect 10968 43726 11020 43732
rect 10048 43308 10100 43314
rect 10048 43250 10100 43256
rect 9956 42832 10008 42838
rect 9956 42774 10008 42780
rect 10980 42770 11008 43726
rect 11072 43314 11100 45222
rect 11716 45082 11744 45358
rect 11704 45076 11756 45082
rect 11704 45018 11756 45024
rect 11152 44940 11204 44946
rect 11152 44882 11204 44888
rect 11164 44402 11192 44882
rect 11244 44872 11296 44878
rect 11244 44814 11296 44820
rect 11256 44538 11284 44814
rect 11244 44532 11296 44538
rect 11244 44474 11296 44480
rect 11152 44396 11204 44402
rect 11152 44338 11204 44344
rect 11060 43308 11112 43314
rect 11060 43250 11112 43256
rect 10968 42764 11020 42770
rect 10968 42706 11020 42712
rect 9496 40724 9548 40730
rect 9496 40666 9548 40672
rect 10692 40724 10744 40730
rect 10692 40666 10744 40672
rect 9680 40044 9732 40050
rect 9680 39986 9732 39992
rect 9692 39642 9720 39986
rect 9680 39636 9732 39642
rect 9680 39578 9732 39584
rect 9220 39432 9272 39438
rect 9220 39374 9272 39380
rect 8668 39296 8720 39302
rect 8668 39238 8720 39244
rect 9036 39296 9088 39302
rect 9036 39238 9088 39244
rect 8680 39030 8708 39238
rect 8208 39024 8260 39030
rect 8208 38966 8260 38972
rect 8668 39024 8720 39030
rect 8668 38966 8720 38972
rect 9048 38962 9076 39238
rect 7472 38956 7524 38962
rect 7472 38898 7524 38904
rect 7840 38956 7892 38962
rect 7840 38898 7892 38904
rect 8024 38956 8076 38962
rect 8024 38898 8076 38904
rect 9036 38956 9088 38962
rect 9036 38898 9088 38904
rect 7288 38344 7340 38350
rect 7288 38286 7340 38292
rect 5448 37936 5500 37942
rect 5448 37878 5500 37884
rect 1676 37868 1728 37874
rect 1676 37810 1728 37816
rect 5356 37800 5408 37806
rect 5356 37742 5408 37748
rect 4804 37664 4856 37670
rect 4804 37606 4856 37612
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4816 36786 4844 37606
rect 5264 37188 5316 37194
rect 5264 37130 5316 37136
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 5276 36922 5304 37130
rect 5264 36916 5316 36922
rect 5264 36858 5316 36864
rect 5368 36802 5396 37742
rect 5460 37194 5488 37878
rect 7012 37800 7064 37806
rect 7012 37742 7064 37748
rect 5632 37664 5684 37670
rect 5632 37606 5684 37612
rect 5448 37188 5500 37194
rect 5448 37130 5500 37136
rect 4804 36780 4856 36786
rect 4804 36722 4856 36728
rect 5276 36774 5396 36802
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4804 36032 4856 36038
rect 4804 35974 4856 35980
rect 4816 35714 4844 35974
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 5276 35894 5304 36774
rect 5460 36258 5488 37130
rect 5644 36786 5672 37606
rect 7024 37262 7052 37742
rect 7300 37738 7328 38286
rect 8036 37806 8064 38898
rect 9048 38554 9076 38898
rect 9232 38554 9260 39374
rect 10704 39370 10732 40666
rect 10876 40656 10928 40662
rect 10876 40598 10928 40604
rect 10888 39506 10916 40598
rect 10968 40520 11020 40526
rect 10968 40462 11020 40468
rect 10980 40186 11008 40462
rect 10968 40180 11020 40186
rect 10968 40122 11020 40128
rect 11164 40066 11192 44338
rect 11716 44334 11744 45018
rect 11808 44538 11836 45426
rect 11900 44878 11928 45426
rect 13820 45280 13872 45286
rect 13820 45222 13872 45228
rect 11888 44872 11940 44878
rect 11888 44814 11940 44820
rect 11796 44532 11848 44538
rect 11796 44474 11848 44480
rect 11704 44328 11756 44334
rect 11704 44270 11756 44276
rect 11520 44260 11572 44266
rect 11520 44202 11572 44208
rect 11336 42764 11388 42770
rect 11336 42706 11388 42712
rect 11348 42634 11376 42706
rect 11336 42628 11388 42634
rect 11336 42570 11388 42576
rect 11532 41414 11560 44202
rect 11612 43648 11664 43654
rect 11612 43590 11664 43596
rect 11624 43314 11652 43590
rect 11612 43308 11664 43314
rect 11612 43250 11664 43256
rect 11716 42906 11744 44270
rect 11808 44198 11836 44474
rect 11900 44334 11928 44814
rect 12532 44804 12584 44810
rect 12532 44746 12584 44752
rect 12256 44736 12308 44742
rect 12256 44678 12308 44684
rect 12440 44736 12492 44742
rect 12440 44678 12492 44684
rect 11888 44328 11940 44334
rect 11888 44270 11940 44276
rect 11796 44192 11848 44198
rect 11796 44134 11848 44140
rect 11808 43994 11836 44134
rect 11796 43988 11848 43994
rect 11796 43930 11848 43936
rect 12268 43790 12296 44678
rect 12452 44470 12480 44678
rect 12440 44464 12492 44470
rect 12440 44406 12492 44412
rect 12544 43926 12572 44746
rect 13832 44470 13860 45222
rect 13820 44464 13872 44470
rect 13820 44406 13872 44412
rect 12716 44396 12768 44402
rect 12716 44338 12768 44344
rect 13452 44396 13504 44402
rect 13452 44338 13504 44344
rect 12728 43926 12756 44338
rect 12900 44192 12952 44198
rect 12900 44134 12952 44140
rect 12912 43994 12940 44134
rect 13464 44010 13492 44338
rect 13372 43994 13492 44010
rect 12900 43988 12952 43994
rect 12900 43930 12952 43936
rect 13360 43988 13492 43994
rect 13412 43982 13492 43988
rect 13360 43930 13412 43936
rect 12532 43920 12584 43926
rect 12532 43862 12584 43868
rect 12716 43920 12768 43926
rect 12716 43862 12768 43868
rect 13176 43920 13228 43926
rect 13176 43862 13228 43868
rect 11796 43784 11848 43790
rect 11796 43726 11848 43732
rect 11888 43784 11940 43790
rect 11888 43726 11940 43732
rect 11980 43784 12032 43790
rect 11980 43726 12032 43732
rect 12256 43784 12308 43790
rect 12256 43726 12308 43732
rect 11808 43110 11836 43726
rect 11900 43382 11928 43726
rect 11992 43450 12020 43726
rect 11980 43444 12032 43450
rect 11980 43386 12032 43392
rect 11888 43376 11940 43382
rect 11888 43318 11940 43324
rect 11980 43172 12032 43178
rect 11980 43114 12032 43120
rect 11796 43104 11848 43110
rect 11796 43046 11848 43052
rect 11704 42900 11756 42906
rect 11704 42842 11756 42848
rect 11808 42702 11836 43046
rect 11992 42702 12020 43114
rect 12072 42764 12124 42770
rect 12072 42706 12124 42712
rect 11796 42696 11848 42702
rect 11796 42638 11848 42644
rect 11980 42696 12032 42702
rect 11980 42638 12032 42644
rect 11532 41386 11652 41414
rect 11624 40186 11652 41386
rect 11612 40180 11664 40186
rect 11612 40122 11664 40128
rect 11072 40038 11192 40066
rect 11244 40044 11296 40050
rect 10876 39500 10928 39506
rect 10876 39442 10928 39448
rect 10784 39432 10836 39438
rect 10784 39374 10836 39380
rect 10692 39364 10744 39370
rect 10692 39306 10744 39312
rect 10796 39098 10824 39374
rect 10784 39092 10836 39098
rect 10784 39034 10836 39040
rect 11072 38962 11100 40038
rect 11244 39986 11296 39992
rect 11152 39908 11204 39914
rect 11152 39850 11204 39856
rect 10508 38956 10560 38962
rect 10508 38898 10560 38904
rect 11060 38956 11112 38962
rect 11060 38898 11112 38904
rect 10048 38752 10100 38758
rect 10048 38694 10100 38700
rect 9036 38548 9088 38554
rect 9036 38490 9088 38496
rect 9220 38548 9272 38554
rect 9220 38490 9272 38496
rect 9588 38548 9640 38554
rect 9588 38490 9640 38496
rect 9048 38010 9076 38490
rect 9036 38004 9088 38010
rect 9036 37946 9088 37952
rect 9600 37942 9628 38490
rect 10060 38418 10088 38694
rect 10048 38412 10100 38418
rect 10048 38354 10100 38360
rect 10520 38350 10548 38898
rect 10600 38888 10652 38894
rect 10600 38830 10652 38836
rect 10508 38344 10560 38350
rect 10508 38286 10560 38292
rect 10324 38208 10376 38214
rect 10324 38150 10376 38156
rect 9588 37936 9640 37942
rect 9588 37878 9640 37884
rect 9036 37868 9088 37874
rect 9036 37810 9088 37816
rect 8024 37800 8076 37806
rect 8024 37742 8076 37748
rect 7288 37732 7340 37738
rect 7288 37674 7340 37680
rect 7012 37256 7064 37262
rect 7012 37198 7064 37204
rect 6368 37120 6420 37126
rect 6368 37062 6420 37068
rect 5632 36780 5684 36786
rect 5632 36722 5684 36728
rect 6380 36718 6408 37062
rect 6368 36712 6420 36718
rect 6368 36654 6420 36660
rect 5632 36576 5684 36582
rect 5632 36518 5684 36524
rect 5368 36230 5488 36258
rect 5368 36174 5396 36230
rect 5356 36168 5408 36174
rect 5356 36110 5408 36116
rect 5540 36100 5592 36106
rect 5540 36042 5592 36048
rect 5276 35866 5396 35894
rect 4816 35698 5028 35714
rect 4804 35692 5040 35698
rect 4856 35686 4988 35692
rect 4804 35634 4856 35640
rect 4988 35634 5040 35640
rect 5264 35488 5316 35494
rect 5264 35430 5316 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 5276 34610 5304 35430
rect 5368 35290 5396 35866
rect 5552 35834 5580 36042
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5644 35766 5672 36518
rect 6092 36032 6144 36038
rect 6092 35974 6144 35980
rect 5632 35760 5684 35766
rect 5632 35702 5684 35708
rect 5540 35692 5592 35698
rect 5540 35634 5592 35640
rect 5552 35578 5580 35634
rect 6104 35630 6132 35974
rect 6092 35624 6144 35630
rect 5552 35550 5672 35578
rect 6092 35566 6144 35572
rect 5540 35488 5592 35494
rect 5540 35430 5592 35436
rect 5356 35284 5408 35290
rect 5356 35226 5408 35232
rect 5552 35154 5580 35430
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 5448 34944 5500 34950
rect 5448 34886 5500 34892
rect 5264 34604 5316 34610
rect 5264 34546 5316 34552
rect 4896 34400 4948 34406
rect 4896 34342 4948 34348
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4908 33930 4936 34342
rect 4896 33924 4948 33930
rect 4896 33866 4948 33872
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 5460 32910 5488 34886
rect 5644 34728 5672 35550
rect 6104 35494 6132 35566
rect 6092 35488 6144 35494
rect 6092 35430 6144 35436
rect 6380 35222 6408 36654
rect 6460 36168 6512 36174
rect 6460 36110 6512 36116
rect 6472 35834 6500 36110
rect 6920 36032 6972 36038
rect 6920 35974 6972 35980
rect 6460 35828 6512 35834
rect 6460 35770 6512 35776
rect 6368 35216 6420 35222
rect 6368 35158 6420 35164
rect 5816 35012 5868 35018
rect 5816 34954 5868 34960
rect 5908 35012 5960 35018
rect 5908 34954 5960 34960
rect 5724 34740 5776 34746
rect 5644 34700 5724 34728
rect 5724 34682 5776 34688
rect 5632 34604 5684 34610
rect 5632 34546 5684 34552
rect 5644 34202 5672 34546
rect 5736 34542 5764 34682
rect 5724 34536 5776 34542
rect 5724 34478 5776 34484
rect 5632 34196 5684 34202
rect 5632 34138 5684 34144
rect 5644 33522 5672 34138
rect 5632 33516 5684 33522
rect 5632 33458 5684 33464
rect 5540 33312 5592 33318
rect 5540 33254 5592 33260
rect 5448 32904 5500 32910
rect 5448 32846 5500 32852
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 5552 32434 5580 33254
rect 5644 32910 5672 33458
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5736 32434 5764 34478
rect 5828 34202 5856 34954
rect 5816 34196 5868 34202
rect 5816 34138 5868 34144
rect 5540 32428 5592 32434
rect 5540 32370 5592 32376
rect 5724 32428 5776 32434
rect 5724 32370 5776 32376
rect 848 32224 900 32230
rect 846 32192 848 32201
rect 5632 32224 5684 32230
rect 900 32192 902 32201
rect 5632 32166 5684 32172
rect 846 32127 902 32136
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 5644 31754 5672 32166
rect 5920 32042 5948 34954
rect 6472 34950 6500 35770
rect 6932 35766 6960 35974
rect 6920 35760 6972 35766
rect 6920 35702 6972 35708
rect 8036 35698 8064 37742
rect 9048 37330 9076 37810
rect 9036 37324 9088 37330
rect 9036 37266 9088 37272
rect 8024 35692 8076 35698
rect 8024 35634 8076 35640
rect 6552 35624 6604 35630
rect 6552 35566 6604 35572
rect 6564 34950 6592 35566
rect 6920 35488 6972 35494
rect 6920 35430 6972 35436
rect 6828 35216 6880 35222
rect 6828 35158 6880 35164
rect 6184 34944 6236 34950
rect 6184 34886 6236 34892
rect 6460 34944 6512 34950
rect 6460 34886 6512 34892
rect 6552 34944 6604 34950
rect 6552 34886 6604 34892
rect 6196 34678 6224 34886
rect 6184 34672 6236 34678
rect 6184 34614 6236 34620
rect 6472 34542 6500 34886
rect 6840 34746 6868 35158
rect 6932 34950 6960 35430
rect 7012 35080 7064 35086
rect 7012 35022 7064 35028
rect 6920 34944 6972 34950
rect 6920 34886 6972 34892
rect 7024 34746 7052 35022
rect 6828 34740 6880 34746
rect 6828 34682 6880 34688
rect 7012 34740 7064 34746
rect 7012 34682 7064 34688
rect 6736 34604 6788 34610
rect 6736 34546 6788 34552
rect 6828 34604 6880 34610
rect 6828 34546 6880 34552
rect 6460 34536 6512 34542
rect 6460 34478 6512 34484
rect 6748 33046 6776 34546
rect 6736 33040 6788 33046
rect 6736 32982 6788 32988
rect 6840 32978 6868 34546
rect 9048 34474 9076 37266
rect 10336 37262 10364 38150
rect 10520 38010 10548 38286
rect 10508 38004 10560 38010
rect 10508 37946 10560 37952
rect 10508 37664 10560 37670
rect 10508 37606 10560 37612
rect 10324 37256 10376 37262
rect 10324 37198 10376 37204
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9128 35012 9180 35018
rect 9128 34954 9180 34960
rect 9036 34468 9088 34474
rect 9036 34410 9088 34416
rect 7932 34400 7984 34406
rect 7932 34342 7984 34348
rect 6920 33992 6972 33998
rect 6920 33934 6972 33940
rect 7196 33992 7248 33998
rect 7196 33934 7248 33940
rect 6932 33114 6960 33934
rect 7208 33318 7236 33934
rect 7944 33930 7972 34342
rect 7932 33924 7984 33930
rect 7932 33866 7984 33872
rect 9048 33658 9076 34410
rect 9140 33998 9168 34954
rect 9416 34542 9444 35022
rect 10520 34678 10548 37606
rect 10612 34746 10640 38830
rect 11060 38480 11112 38486
rect 11060 38422 11112 38428
rect 11072 37330 11100 38422
rect 11164 37874 11192 39850
rect 11256 37874 11284 39986
rect 11428 39976 11480 39982
rect 11428 39918 11480 39924
rect 11440 39506 11468 39918
rect 12084 39506 12112 42706
rect 11428 39500 11480 39506
rect 11428 39442 11480 39448
rect 12072 39500 12124 39506
rect 12072 39442 12124 39448
rect 11152 37868 11204 37874
rect 11152 37810 11204 37816
rect 11244 37868 11296 37874
rect 11244 37810 11296 37816
rect 11164 37466 11192 37810
rect 11152 37460 11204 37466
rect 11152 37402 11204 37408
rect 11060 37324 11112 37330
rect 11060 37266 11112 37272
rect 11256 36786 11284 37810
rect 11440 37398 11468 39442
rect 12084 38962 12112 39442
rect 12072 38956 12124 38962
rect 12072 38898 12124 38904
rect 11888 38888 11940 38894
rect 11888 38830 11940 38836
rect 11796 38752 11848 38758
rect 11796 38694 11848 38700
rect 11808 37874 11836 38694
rect 11900 37874 11928 38830
rect 12164 38752 12216 38758
rect 12164 38694 12216 38700
rect 12176 38350 12204 38694
rect 12164 38344 12216 38350
rect 12164 38286 12216 38292
rect 12268 38214 12296 43726
rect 12544 43314 12572 43862
rect 13188 43450 13216 43862
rect 13832 43858 13860 44406
rect 13820 43852 13872 43858
rect 13820 43794 13872 43800
rect 13544 43784 13596 43790
rect 13544 43726 13596 43732
rect 13176 43444 13228 43450
rect 13176 43386 13228 43392
rect 13556 43314 13584 43726
rect 13924 43382 13952 45426
rect 14372 45416 14424 45422
rect 14372 45358 14424 45364
rect 14096 45348 14148 45354
rect 14096 45290 14148 45296
rect 14108 44538 14136 45290
rect 14280 44804 14332 44810
rect 14280 44746 14332 44752
rect 14096 44532 14148 44538
rect 14096 44474 14148 44480
rect 14292 44402 14320 44746
rect 14280 44396 14332 44402
rect 14280 44338 14332 44344
rect 14004 44192 14056 44198
rect 14004 44134 14056 44140
rect 13912 43376 13964 43382
rect 13912 43318 13964 43324
rect 14016 43314 14044 44134
rect 14384 43858 14412 45358
rect 14648 45280 14700 45286
rect 14648 45222 14700 45228
rect 14660 44810 14688 45222
rect 14648 44804 14700 44810
rect 14648 44746 14700 44752
rect 14752 44538 14780 45426
rect 15752 45416 15804 45422
rect 15752 45358 15804 45364
rect 14924 45280 14976 45286
rect 14924 45222 14976 45228
rect 14740 44532 14792 44538
rect 14740 44474 14792 44480
rect 14740 44260 14792 44266
rect 14740 44202 14792 44208
rect 14752 43926 14780 44202
rect 14740 43920 14792 43926
rect 14740 43862 14792 43868
rect 14096 43852 14148 43858
rect 14096 43794 14148 43800
rect 14372 43852 14424 43858
rect 14372 43794 14424 43800
rect 12532 43308 12584 43314
rect 12532 43250 12584 43256
rect 13544 43308 13596 43314
rect 13544 43250 13596 43256
rect 14004 43308 14056 43314
rect 14004 43250 14056 43256
rect 12624 43240 12676 43246
rect 12624 43182 12676 43188
rect 12440 43104 12492 43110
rect 12440 43046 12492 43052
rect 12452 42702 12480 43046
rect 12440 42696 12492 42702
rect 12440 42638 12492 42644
rect 12636 41614 12664 43182
rect 13556 42702 13584 43250
rect 14108 43246 14136 43794
rect 14096 43240 14148 43246
rect 14096 43182 14148 43188
rect 14648 43172 14700 43178
rect 14648 43114 14700 43120
rect 14660 42702 14688 43114
rect 13544 42696 13596 42702
rect 13544 42638 13596 42644
rect 14096 42696 14148 42702
rect 14096 42638 14148 42644
rect 14648 42696 14700 42702
rect 14648 42638 14700 42644
rect 12624 41608 12676 41614
rect 12624 41550 12676 41556
rect 13176 39976 13228 39982
rect 13176 39918 13228 39924
rect 13188 39098 13216 39918
rect 13636 39432 13688 39438
rect 13636 39374 13688 39380
rect 13176 39092 13228 39098
rect 13176 39034 13228 39040
rect 13648 38962 13676 39374
rect 14108 38962 14136 42638
rect 14752 42566 14780 43862
rect 14936 42888 14964 45222
rect 15016 44872 15068 44878
rect 15016 44814 15068 44820
rect 15028 43858 15056 44814
rect 15764 44402 15792 45358
rect 16040 45082 16068 45426
rect 18144 45416 18196 45422
rect 18144 45358 18196 45364
rect 18420 45416 18472 45422
rect 18420 45358 18472 45364
rect 16488 45280 16540 45286
rect 16488 45222 16540 45228
rect 17500 45280 17552 45286
rect 17500 45222 17552 45228
rect 17776 45280 17828 45286
rect 17776 45222 17828 45228
rect 16028 45076 16080 45082
rect 16028 45018 16080 45024
rect 16500 44470 16528 45222
rect 17512 44810 17540 45222
rect 17500 44804 17552 44810
rect 17500 44746 17552 44752
rect 17788 44538 17816 45222
rect 18156 44742 18184 45358
rect 18432 44878 18460 45358
rect 18420 44872 18472 44878
rect 18420 44814 18472 44820
rect 19340 44872 19392 44878
rect 19340 44814 19392 44820
rect 18144 44736 18196 44742
rect 18144 44678 18196 44684
rect 17776 44532 17828 44538
rect 17776 44474 17828 44480
rect 16488 44464 16540 44470
rect 16488 44406 16540 44412
rect 15752 44396 15804 44402
rect 15752 44338 15804 44344
rect 15568 44328 15620 44334
rect 15568 44270 15620 44276
rect 15016 43852 15068 43858
rect 15016 43794 15068 43800
rect 15580 43790 15608 44270
rect 15568 43784 15620 43790
rect 15568 43726 15620 43732
rect 15200 43240 15252 43246
rect 15200 43182 15252 43188
rect 14936 42860 15056 42888
rect 15028 42702 15056 42860
rect 15212 42770 15240 43182
rect 15200 42764 15252 42770
rect 15200 42706 15252 42712
rect 15016 42696 15068 42702
rect 15016 42638 15068 42644
rect 15580 42634 15608 43726
rect 15568 42628 15620 42634
rect 15568 42570 15620 42576
rect 14740 42560 14792 42566
rect 14740 42502 14792 42508
rect 15580 40050 15608 42570
rect 15292 40044 15344 40050
rect 15292 39986 15344 39992
rect 15568 40044 15620 40050
rect 15568 39986 15620 39992
rect 15200 39976 15252 39982
rect 15200 39918 15252 39924
rect 15212 39370 15240 39918
rect 15304 39574 15332 39986
rect 15764 39914 15792 44338
rect 15844 43716 15896 43722
rect 15844 43658 15896 43664
rect 15856 43450 15884 43658
rect 16500 43654 16528 44406
rect 18052 44396 18104 44402
rect 18052 44338 18104 44344
rect 16856 44328 16908 44334
rect 16856 44270 16908 44276
rect 16672 43784 16724 43790
rect 16672 43726 16724 43732
rect 16764 43784 16816 43790
rect 16764 43726 16816 43732
rect 16396 43648 16448 43654
rect 16396 43590 16448 43596
rect 16488 43648 16540 43654
rect 16488 43590 16540 43596
rect 15844 43444 15896 43450
rect 15844 43386 15896 43392
rect 16120 42696 16172 42702
rect 16120 42638 16172 42644
rect 16028 41472 16080 41478
rect 16028 41414 16080 41420
rect 16040 40526 16068 41414
rect 16028 40520 16080 40526
rect 16028 40462 16080 40468
rect 15844 40452 15896 40458
rect 15844 40394 15896 40400
rect 15752 39908 15804 39914
rect 15752 39850 15804 39856
rect 15660 39840 15712 39846
rect 15660 39782 15712 39788
rect 15292 39568 15344 39574
rect 15292 39510 15344 39516
rect 15200 39364 15252 39370
rect 15200 39306 15252 39312
rect 12716 38956 12768 38962
rect 12716 38898 12768 38904
rect 13636 38956 13688 38962
rect 13636 38898 13688 38904
rect 13912 38956 13964 38962
rect 13912 38898 13964 38904
rect 14096 38956 14148 38962
rect 14096 38898 14148 38904
rect 12532 38820 12584 38826
rect 12532 38762 12584 38768
rect 12348 38752 12400 38758
rect 12348 38694 12400 38700
rect 12360 38282 12388 38694
rect 12348 38276 12400 38282
rect 12348 38218 12400 38224
rect 12256 38208 12308 38214
rect 12256 38150 12308 38156
rect 12360 37874 12388 38218
rect 11796 37868 11848 37874
rect 11796 37810 11848 37816
rect 11888 37868 11940 37874
rect 11888 37810 11940 37816
rect 12348 37868 12400 37874
rect 12348 37810 12400 37816
rect 11428 37392 11480 37398
rect 11428 37334 11480 37340
rect 12360 37330 12388 37810
rect 12440 37460 12492 37466
rect 12440 37402 12492 37408
rect 12348 37324 12400 37330
rect 12348 37266 12400 37272
rect 12360 36854 12388 37266
rect 12348 36848 12400 36854
rect 12348 36790 12400 36796
rect 12452 36786 12480 37402
rect 11244 36780 11296 36786
rect 11244 36722 11296 36728
rect 11704 36780 11756 36786
rect 11704 36722 11756 36728
rect 12440 36780 12492 36786
rect 12440 36722 12492 36728
rect 11716 35290 11744 36722
rect 12544 36650 12572 38762
rect 12728 38554 12756 38898
rect 12808 38888 12860 38894
rect 12808 38830 12860 38836
rect 13176 38888 13228 38894
rect 13176 38830 13228 38836
rect 12716 38548 12768 38554
rect 12716 38490 12768 38496
rect 12624 37800 12676 37806
rect 12624 37742 12676 37748
rect 12532 36644 12584 36650
rect 12532 36586 12584 36592
rect 11704 35284 11756 35290
rect 11704 35226 11756 35232
rect 11888 35080 11940 35086
rect 11888 35022 11940 35028
rect 12072 35080 12124 35086
rect 12072 35022 12124 35028
rect 10600 34740 10652 34746
rect 10600 34682 10652 34688
rect 10508 34672 10560 34678
rect 10508 34614 10560 34620
rect 10876 34672 10928 34678
rect 10876 34614 10928 34620
rect 9864 34604 9916 34610
rect 9864 34546 9916 34552
rect 10140 34604 10192 34610
rect 10140 34546 10192 34552
rect 10784 34604 10836 34610
rect 10784 34546 10836 34552
rect 9404 34536 9456 34542
rect 9404 34478 9456 34484
rect 9680 34536 9732 34542
rect 9680 34478 9732 34484
rect 9128 33992 9180 33998
rect 9128 33934 9180 33940
rect 9036 33652 9088 33658
rect 9036 33594 9088 33600
rect 7196 33312 7248 33318
rect 7196 33254 7248 33260
rect 6920 33108 6972 33114
rect 6920 33050 6972 33056
rect 6828 32972 6880 32978
rect 6828 32914 6880 32920
rect 6460 32904 6512 32910
rect 6460 32846 6512 32852
rect 6472 32570 6500 32846
rect 6460 32564 6512 32570
rect 6460 32506 6512 32512
rect 6644 32428 6696 32434
rect 6644 32370 6696 32376
rect 5920 32026 6040 32042
rect 5920 32020 6052 32026
rect 5920 32014 6000 32020
rect 5632 31748 5684 31754
rect 5632 31690 5684 31696
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 5920 31346 5948 32014
rect 6000 31962 6052 31968
rect 6656 31754 6684 32370
rect 6644 31748 6696 31754
rect 6644 31690 6696 31696
rect 6656 31346 6684 31690
rect 6840 31346 6868 32914
rect 7208 32842 7236 33254
rect 9416 32910 9444 34478
rect 9692 34202 9720 34478
rect 9680 34196 9732 34202
rect 9680 34138 9732 34144
rect 9692 33522 9720 34138
rect 9876 33522 9904 34546
rect 9956 34536 10008 34542
rect 9956 34478 10008 34484
rect 9968 34202 9996 34478
rect 9956 34196 10008 34202
rect 9956 34138 10008 34144
rect 9968 33658 9996 34138
rect 9956 33652 10008 33658
rect 9956 33594 10008 33600
rect 9680 33516 9732 33522
rect 9680 33458 9732 33464
rect 9864 33516 9916 33522
rect 9864 33458 9916 33464
rect 9876 32978 9904 33458
rect 9968 32978 9996 33594
rect 10152 33590 10180 34546
rect 10692 33992 10744 33998
rect 10692 33934 10744 33940
rect 10140 33584 10192 33590
rect 10140 33526 10192 33532
rect 9864 32972 9916 32978
rect 9864 32914 9916 32920
rect 9956 32972 10008 32978
rect 9956 32914 10008 32920
rect 9404 32904 9456 32910
rect 9404 32846 9456 32852
rect 7196 32836 7248 32842
rect 7196 32778 7248 32784
rect 7208 32230 7236 32778
rect 10152 32502 10180 33526
rect 10600 33448 10652 33454
rect 10600 33390 10652 33396
rect 10612 32570 10640 33390
rect 10704 33046 10732 33934
rect 10796 33114 10824 34546
rect 10784 33108 10836 33114
rect 10784 33050 10836 33056
rect 10692 33040 10744 33046
rect 10692 32982 10744 32988
rect 10600 32564 10652 32570
rect 10600 32506 10652 32512
rect 10796 32502 10824 33050
rect 10140 32496 10192 32502
rect 10140 32438 10192 32444
rect 10784 32496 10836 32502
rect 10784 32438 10836 32444
rect 10888 32434 10916 34614
rect 11244 34536 11296 34542
rect 11244 34478 11296 34484
rect 11256 33998 11284 34478
rect 11244 33992 11296 33998
rect 11244 33934 11296 33940
rect 11520 33992 11572 33998
rect 11520 33934 11572 33940
rect 11532 33658 11560 33934
rect 11520 33652 11572 33658
rect 11520 33594 11572 33600
rect 11900 33590 11928 35022
rect 11704 33584 11756 33590
rect 11704 33526 11756 33532
rect 11888 33584 11940 33590
rect 11888 33526 11940 33532
rect 11060 33312 11112 33318
rect 11060 33254 11112 33260
rect 7932 32428 7984 32434
rect 7932 32370 7984 32376
rect 10876 32428 10928 32434
rect 10876 32370 10928 32376
rect 7196 32224 7248 32230
rect 7196 32166 7248 32172
rect 7208 31822 7236 32166
rect 7944 32026 7972 32370
rect 11072 32298 11100 33254
rect 11716 32570 11744 33526
rect 12084 33386 12112 35022
rect 12348 34944 12400 34950
rect 12348 34886 12400 34892
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 12072 33380 12124 33386
rect 12072 33322 12124 33328
rect 11888 33312 11940 33318
rect 11888 33254 11940 33260
rect 11900 32978 11928 33254
rect 11888 32972 11940 32978
rect 11888 32914 11940 32920
rect 12084 32570 12112 33322
rect 12164 32768 12216 32774
rect 12164 32710 12216 32716
rect 11704 32564 11756 32570
rect 11704 32506 11756 32512
rect 12072 32564 12124 32570
rect 12072 32506 12124 32512
rect 11060 32292 11112 32298
rect 11060 32234 11112 32240
rect 7932 32020 7984 32026
rect 7932 31962 7984 31968
rect 12176 31822 12204 32710
rect 12268 32230 12296 34546
rect 12360 34202 12388 34886
rect 12348 34196 12400 34202
rect 12348 34138 12400 34144
rect 12360 33114 12388 34138
rect 12636 34134 12664 37742
rect 12728 37312 12756 38490
rect 12820 38010 12848 38830
rect 13188 38350 13216 38830
rect 12900 38344 12952 38350
rect 12900 38286 12952 38292
rect 13084 38344 13136 38350
rect 13084 38286 13136 38292
rect 13176 38344 13228 38350
rect 13176 38286 13228 38292
rect 12808 38004 12860 38010
rect 12808 37946 12860 37952
rect 12912 37466 12940 38286
rect 13096 38010 13124 38286
rect 13084 38004 13136 38010
rect 13084 37946 13136 37952
rect 12992 37936 13044 37942
rect 12992 37878 13044 37884
rect 12900 37460 12952 37466
rect 12900 37402 12952 37408
rect 12808 37324 12860 37330
rect 12728 37284 12808 37312
rect 12808 37266 12860 37272
rect 12820 34678 12848 37266
rect 12900 37256 12952 37262
rect 12900 37198 12952 37204
rect 12912 36922 12940 37198
rect 12900 36916 12952 36922
rect 12900 36858 12952 36864
rect 13004 35154 13032 37878
rect 13924 37398 13952 38898
rect 14004 38752 14056 38758
rect 14004 38694 14056 38700
rect 14016 38350 14044 38694
rect 14004 38344 14056 38350
rect 14004 38286 14056 38292
rect 14108 38010 14136 38898
rect 15304 38418 15332 39510
rect 15672 39438 15700 39782
rect 15856 39438 15884 40394
rect 15476 39432 15528 39438
rect 15476 39374 15528 39380
rect 15660 39432 15712 39438
rect 15660 39374 15712 39380
rect 15844 39432 15896 39438
rect 15844 39374 15896 39380
rect 15384 38752 15436 38758
rect 15384 38694 15436 38700
rect 15292 38412 15344 38418
rect 15292 38354 15344 38360
rect 14096 38004 14148 38010
rect 14096 37946 14148 37952
rect 13912 37392 13964 37398
rect 13912 37334 13964 37340
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 12992 35148 13044 35154
rect 12992 35090 13044 35096
rect 13004 34746 13032 35090
rect 12992 34740 13044 34746
rect 12992 34682 13044 34688
rect 12808 34672 12860 34678
rect 12808 34614 12860 34620
rect 12624 34128 12676 34134
rect 12624 34070 12676 34076
rect 13004 33998 13032 34682
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12716 33992 12768 33998
rect 12716 33934 12768 33940
rect 12992 33992 13044 33998
rect 12992 33934 13044 33940
rect 12440 33856 12492 33862
rect 12440 33798 12492 33804
rect 12452 33522 12480 33798
rect 12440 33516 12492 33522
rect 12440 33458 12492 33464
rect 12544 33386 12572 33934
rect 12532 33380 12584 33386
rect 12532 33322 12584 33328
rect 12348 33108 12400 33114
rect 12348 33050 12400 33056
rect 12360 32910 12388 33050
rect 12348 32904 12400 32910
rect 12348 32846 12400 32852
rect 12544 32570 12572 33322
rect 12532 32564 12584 32570
rect 12532 32506 12584 32512
rect 12256 32224 12308 32230
rect 12256 32166 12308 32172
rect 12728 32026 12756 33934
rect 12808 33924 12860 33930
rect 12808 33866 12860 33872
rect 12716 32020 12768 32026
rect 12716 31962 12768 31968
rect 12820 31822 12848 33866
rect 7196 31816 7248 31822
rect 7196 31758 7248 31764
rect 8300 31816 8352 31822
rect 8300 31758 8352 31764
rect 12164 31816 12216 31822
rect 12164 31758 12216 31764
rect 12808 31816 12860 31822
rect 12808 31758 12860 31764
rect 5908 31340 5960 31346
rect 5908 31282 5960 31288
rect 6644 31340 6696 31346
rect 6644 31282 6696 31288
rect 6828 31340 6880 31346
rect 6828 31282 6880 31288
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 6656 30598 6684 31282
rect 6840 31226 6868 31282
rect 6748 31198 6868 31226
rect 6748 30938 6776 31198
rect 6828 31136 6880 31142
rect 6828 31078 6880 31084
rect 6736 30932 6788 30938
rect 6736 30874 6788 30880
rect 6840 30734 6868 31078
rect 7208 30734 7236 31758
rect 8312 31482 8340 31758
rect 8300 31476 8352 31482
rect 8300 31418 8352 31424
rect 6828 30728 6880 30734
rect 6828 30670 6880 30676
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 6644 30592 6696 30598
rect 6644 30534 6696 30540
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 1308 30252 1360 30258
rect 1308 30194 1360 30200
rect 1320 30025 1348 30194
rect 1676 30048 1728 30054
rect 1306 30016 1362 30025
rect 1676 29990 1728 29996
rect 1306 29951 1362 29960
rect 848 29640 900 29646
rect 848 29582 900 29588
rect 860 29481 888 29582
rect 846 29472 902 29481
rect 846 29407 902 29416
rect 1688 29170 1716 29990
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 1676 29164 1728 29170
rect 1676 29106 1728 29112
rect 4804 29028 4856 29034
rect 4804 28970 4856 28976
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4816 28490 4844 28970
rect 7208 28490 7236 30670
rect 8484 30592 8536 30598
rect 8484 30534 8536 30540
rect 8496 30054 8524 30534
rect 9036 30184 9088 30190
rect 9036 30126 9088 30132
rect 8484 30048 8536 30054
rect 8484 29990 8536 29996
rect 8496 29646 8524 29990
rect 9048 29782 9076 30126
rect 9404 30048 9456 30054
rect 9404 29990 9456 29996
rect 9036 29776 9088 29782
rect 9036 29718 9088 29724
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 8300 29232 8352 29238
rect 8300 29174 8352 29180
rect 8312 28558 8340 29174
rect 8496 29170 8524 29582
rect 8484 29164 8536 29170
rect 8484 29106 8536 29112
rect 9048 28642 9076 29718
rect 9048 28614 9168 28642
rect 9416 28626 9444 29990
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 10324 29640 10376 29646
rect 10324 29582 10376 29588
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 9784 28626 9812 29242
rect 10048 29028 10100 29034
rect 10048 28970 10100 28976
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9876 28626 9904 28902
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 4804 28484 4856 28490
rect 4804 28426 4856 28432
rect 7196 28484 7248 28490
rect 7196 28426 7248 28432
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 6840 28082 6868 28358
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 7208 28014 7236 28426
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 8208 28416 8260 28422
rect 8208 28358 8260 28364
rect 7484 28082 7512 28358
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 112 27940 164 27946
rect 112 27882 164 27888
rect 6736 27872 6788 27878
rect 6736 27814 6788 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 6748 27402 6776 27814
rect 7208 27470 7236 27950
rect 8220 27470 8248 28358
rect 8312 27606 8340 28494
rect 9140 28490 9168 28614
rect 9404 28620 9456 28626
rect 9404 28562 9456 28568
rect 9772 28620 9824 28626
rect 9772 28562 9824 28568
rect 9864 28620 9916 28626
rect 9864 28562 9916 28568
rect 8668 28484 8720 28490
rect 8668 28426 8720 28432
rect 9128 28484 9180 28490
rect 9128 28426 9180 28432
rect 8484 28416 8536 28422
rect 8484 28358 8536 28364
rect 8496 28218 8524 28358
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 8300 27600 8352 27606
rect 8300 27542 8352 27548
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 7196 27464 7248 27470
rect 7196 27406 7248 27412
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 6736 27396 6788 27402
rect 6736 27338 6788 27344
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 7208 27062 7236 27406
rect 8404 27130 8432 27474
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 7196 27056 7248 27062
rect 8496 27010 8524 28154
rect 8680 27946 8708 28426
rect 8668 27940 8720 27946
rect 8668 27882 8720 27888
rect 8852 27872 8904 27878
rect 8852 27814 8904 27820
rect 7196 26998 7248 27004
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8312 26982 8524 27010
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 8128 26586 8156 26930
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 8312 26382 8340 26982
rect 8864 26450 8892 27814
rect 9140 27470 9168 28426
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 9404 28416 9456 28422
rect 9404 28358 9456 28364
rect 9324 27674 9352 28358
rect 9312 27668 9364 27674
rect 9312 27610 9364 27616
rect 9416 27538 9444 28358
rect 9404 27532 9456 27538
rect 9404 27474 9456 27480
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 8944 26988 8996 26994
rect 8944 26930 8996 26936
rect 8852 26444 8904 26450
rect 8852 26386 8904 26392
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 8312 25702 8340 26318
rect 8956 26042 8984 26930
rect 9416 26450 9444 27474
rect 9876 27062 9904 28562
rect 10060 28490 10088 28970
rect 10336 28966 10364 29582
rect 10520 29306 10548 29650
rect 10508 29300 10560 29306
rect 10508 29242 10560 29248
rect 10324 28960 10376 28966
rect 10324 28902 10376 28908
rect 10140 28756 10192 28762
rect 10140 28698 10192 28704
rect 10048 28484 10100 28490
rect 10048 28426 10100 28432
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 9968 28082 9996 28358
rect 10060 28218 10088 28426
rect 10048 28212 10100 28218
rect 10048 28154 10100 28160
rect 10152 28082 10180 28698
rect 10520 28218 10548 29242
rect 10876 29232 10928 29238
rect 10876 29174 10928 29180
rect 12900 29232 12952 29238
rect 12900 29174 12952 29180
rect 10888 28218 10916 29174
rect 11336 29096 11388 29102
rect 11336 29038 11388 29044
rect 10968 28960 11020 28966
rect 10968 28902 11020 28908
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10876 28212 10928 28218
rect 10876 28154 10928 28160
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 10140 28076 10192 28082
rect 10140 28018 10192 28024
rect 10980 28014 11008 28902
rect 11348 28762 11376 29038
rect 11428 28960 11480 28966
rect 11428 28902 11480 28908
rect 11336 28756 11388 28762
rect 11336 28698 11388 28704
rect 11060 28688 11112 28694
rect 11060 28630 11112 28636
rect 11072 28082 11100 28630
rect 11060 28076 11112 28082
rect 11060 28018 11112 28024
rect 11440 28014 11468 28902
rect 12348 28484 12400 28490
rect 12348 28426 12400 28432
rect 12164 28076 12216 28082
rect 12164 28018 12216 28024
rect 10968 28008 11020 28014
rect 10968 27950 11020 27956
rect 11428 28008 11480 28014
rect 11428 27950 11480 27956
rect 10508 27940 10560 27946
rect 10508 27882 10560 27888
rect 10048 27464 10100 27470
rect 10048 27406 10100 27412
rect 10060 27130 10088 27406
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 9864 27056 9916 27062
rect 9864 26998 9916 27004
rect 10520 26994 10548 27882
rect 10876 27872 10928 27878
rect 10876 27814 10928 27820
rect 10692 27328 10744 27334
rect 10692 27270 10744 27276
rect 10704 27062 10732 27270
rect 10692 27056 10744 27062
rect 10692 26998 10744 27004
rect 10888 26994 10916 27814
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11072 27130 11100 27406
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 11440 27062 11468 27950
rect 12176 27674 12204 28018
rect 12360 27878 12388 28426
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12348 27872 12400 27878
rect 12348 27814 12400 27820
rect 12164 27668 12216 27674
rect 12164 27610 12216 27616
rect 12360 27130 12388 27814
rect 12728 27674 12756 28018
rect 12716 27668 12768 27674
rect 12716 27610 12768 27616
rect 12348 27124 12400 27130
rect 12348 27066 12400 27072
rect 11428 27056 11480 27062
rect 11428 26998 11480 27004
rect 12728 26994 12756 27610
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 9404 26444 9456 26450
rect 9404 26386 9456 26392
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 8944 26036 8996 26042
rect 8944 25978 8996 25984
rect 9324 25906 9352 26182
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 8300 25696 8352 25702
rect 8300 25638 8352 25644
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 848 24200 900 24206
rect 848 24142 900 24148
rect 860 24041 888 24142
rect 846 24032 902 24041
rect 846 23967 902 23976
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 9784 23730 9812 25638
rect 12268 24818 12296 26318
rect 12716 26308 12768 26314
rect 12716 26250 12768 26256
rect 12728 26042 12756 26250
rect 12716 26036 12768 26042
rect 12716 25978 12768 25984
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10612 23730 10640 24006
rect 11072 23866 11100 24142
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 11992 23730 12020 24142
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 11980 23724 12032 23730
rect 11980 23666 12032 23672
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 848 23520 900 23526
rect 848 23462 900 23468
rect 860 23361 888 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 846 23352 902 23361
rect 4214 23355 4522 23364
rect 846 23287 902 23296
rect 8496 23186 8524 23598
rect 8484 23180 8536 23186
rect 8484 23122 8536 23128
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4632 22778 4660 22986
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 1216 22024 1268 22030
rect 1216 21966 1268 21972
rect 1228 21865 1256 21966
rect 4632 21894 4660 22578
rect 5632 22568 5684 22574
rect 5632 22510 5684 22516
rect 4620 21888 4672 21894
rect 1214 21856 1270 21865
rect 4620 21830 4672 21836
rect 1214 21791 1270 21800
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 5644 20058 5672 22510
rect 6472 20466 6500 23054
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8404 22642 8432 22918
rect 8496 22658 8524 23122
rect 8772 22778 8800 23666
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8496 22642 8616 22658
rect 9416 22642 9444 23054
rect 10336 23050 10364 23462
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 8392 22636 8444 22642
rect 8496 22636 8628 22642
rect 8496 22630 8576 22636
rect 8392 22578 8444 22584
rect 8576 22578 8628 22584
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9416 21010 9444 22578
rect 9784 22098 9812 22918
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10704 22234 10732 22578
rect 10888 22438 10916 23462
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 10876 22432 10928 22438
rect 10876 22374 10928 22380
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 10888 22030 10916 22374
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10888 21554 10916 21966
rect 11256 21554 11284 22374
rect 11624 21622 11652 22918
rect 11808 22574 11836 23054
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11612 21616 11664 21622
rect 11612 21558 11664 21564
rect 11808 21554 11836 22510
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6564 20058 6592 20402
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 8128 19922 8156 20198
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18766 4660 19246
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 3804 18426 3832 18702
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 848 18080 900 18086
rect 848 18022 900 18028
rect 860 17921 888 18022
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 846 17912 902 17921
rect 4214 17915 4522 17924
rect 846 17847 902 17856
rect 4632 17814 4660 18702
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4620 17808 4672 17814
rect 4620 17750 4672 17756
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 3160 17338 3188 17614
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3436 17202 3464 17478
rect 4632 17270 4660 17478
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 1308 17196 1360 17202
rect 1308 17138 1360 17144
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 1320 17105 1348 17138
rect 1306 17096 1362 17105
rect 1306 17031 1362 17040
rect 4724 16998 4752 18090
rect 4816 17610 4844 18566
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5276 18358 5304 18702
rect 5264 18352 5316 18358
rect 5264 18294 5316 18300
rect 5276 17678 5304 18294
rect 5460 18290 5488 19110
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5552 17338 5580 18634
rect 5920 17542 5948 19314
rect 6748 18630 6776 19722
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7116 18970 7144 19246
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7116 18714 7144 18906
rect 7576 18766 7604 19654
rect 7852 19514 7880 19790
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 9416 19378 9444 20946
rect 10796 20942 10824 21286
rect 11900 21146 11928 21966
rect 11992 21554 12020 23666
rect 12084 23254 12112 23802
rect 12164 23656 12216 23662
rect 12164 23598 12216 23604
rect 12176 23322 12204 23598
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 12084 21350 12112 23190
rect 12164 23044 12216 23050
rect 12164 22986 12216 22992
rect 12176 22778 12204 22986
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12268 22094 12296 24754
rect 12452 24410 12480 24754
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12636 23322 12664 24142
rect 12728 23730 12756 25978
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12728 23118 12756 23666
rect 12808 23248 12860 23254
rect 12808 23190 12860 23196
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12360 22658 12388 22918
rect 12360 22642 12480 22658
rect 12360 22636 12492 22642
rect 12360 22630 12440 22636
rect 12440 22578 12492 22584
rect 12452 22234 12480 22578
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12544 22098 12572 22918
rect 12176 22066 12296 22094
rect 12532 22092 12584 22098
rect 12176 22030 12204 22066
rect 12532 22034 12584 22040
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 12176 21010 12204 21966
rect 12256 21412 12308 21418
rect 12256 21354 12308 21360
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 12268 20466 12296 21354
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12452 20602 12480 20810
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12544 20534 12572 22034
rect 12636 21690 12664 23054
rect 12820 22642 12848 23190
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12912 21554 12940 29174
rect 13004 29170 13032 33934
rect 13084 33312 13136 33318
rect 13084 33254 13136 33260
rect 13096 32434 13124 33254
rect 13084 32428 13136 32434
rect 13084 32370 13136 32376
rect 13556 29238 13584 37198
rect 13820 33856 13872 33862
rect 13820 33798 13872 33804
rect 13832 33454 13860 33798
rect 13820 33448 13872 33454
rect 13820 33390 13872 33396
rect 14108 33386 14136 37946
rect 15396 37942 15424 38694
rect 14740 37936 14792 37942
rect 14740 37878 14792 37884
rect 15384 37936 15436 37942
rect 15384 37878 15436 37884
rect 14188 37868 14240 37874
rect 14188 37810 14240 37816
rect 14464 37868 14516 37874
rect 14464 37810 14516 37816
rect 14200 37466 14228 37810
rect 14188 37460 14240 37466
rect 14188 37402 14240 37408
rect 14476 37194 14504 37810
rect 14752 37262 14780 37878
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 14648 37256 14700 37262
rect 14648 37198 14700 37204
rect 14740 37256 14792 37262
rect 14740 37198 14792 37204
rect 14464 37188 14516 37194
rect 14464 37130 14516 37136
rect 14660 36922 14688 37198
rect 14648 36916 14700 36922
rect 14648 36858 14700 36864
rect 14752 34746 14780 37198
rect 15212 36922 15240 37810
rect 15488 37738 15516 39374
rect 16040 39370 16068 40462
rect 16132 39642 16160 42638
rect 16304 42628 16356 42634
rect 16304 42570 16356 42576
rect 16316 40730 16344 42570
rect 16304 40724 16356 40730
rect 16304 40666 16356 40672
rect 16408 40202 16436 43590
rect 16488 42560 16540 42566
rect 16488 42502 16540 42508
rect 16212 40180 16264 40186
rect 16212 40122 16264 40128
rect 16316 40174 16436 40202
rect 16120 39636 16172 39642
rect 16120 39578 16172 39584
rect 15568 39364 15620 39370
rect 15568 39306 15620 39312
rect 16028 39364 16080 39370
rect 16028 39306 16080 39312
rect 15580 38894 15608 39306
rect 15844 38956 15896 38962
rect 15844 38898 15896 38904
rect 15568 38888 15620 38894
rect 15568 38830 15620 38836
rect 15580 38486 15608 38830
rect 15568 38480 15620 38486
rect 15568 38422 15620 38428
rect 15856 38350 15884 38898
rect 16224 38350 16252 40122
rect 16316 38962 16344 40174
rect 16396 39840 16448 39846
rect 16396 39782 16448 39788
rect 16408 39438 16436 39782
rect 16500 39522 16528 42502
rect 16684 40186 16712 43726
rect 16776 43450 16804 43726
rect 16868 43722 16896 44270
rect 17684 44260 17736 44266
rect 17684 44202 17736 44208
rect 17696 43790 17724 44202
rect 18064 43994 18092 44338
rect 18052 43988 18104 43994
rect 18052 43930 18104 43936
rect 17132 43784 17184 43790
rect 17132 43726 17184 43732
rect 17684 43784 17736 43790
rect 17684 43726 17736 43732
rect 16856 43716 16908 43722
rect 16856 43658 16908 43664
rect 16948 43716 17000 43722
rect 16948 43658 17000 43664
rect 16764 43444 16816 43450
rect 16764 43386 16816 43392
rect 16960 42906 16988 43658
rect 17040 43308 17092 43314
rect 17040 43250 17092 43256
rect 17052 43110 17080 43250
rect 17144 43178 17172 43726
rect 17868 43716 17920 43722
rect 17868 43658 17920 43664
rect 17224 43648 17276 43654
rect 17224 43590 17276 43596
rect 17236 43314 17264 43590
rect 17224 43308 17276 43314
rect 17224 43250 17276 43256
rect 17132 43172 17184 43178
rect 17132 43114 17184 43120
rect 17040 43104 17092 43110
rect 17040 43046 17092 43052
rect 16948 42900 17000 42906
rect 16948 42842 17000 42848
rect 17052 42634 17080 43046
rect 17040 42628 17092 42634
rect 17040 42570 17092 42576
rect 17880 42566 17908 43658
rect 17960 43308 18012 43314
rect 17960 43250 18012 43256
rect 17972 42838 18000 43250
rect 17960 42832 18012 42838
rect 17960 42774 18012 42780
rect 17868 42560 17920 42566
rect 17868 42502 17920 42508
rect 16672 40180 16724 40186
rect 16672 40122 16724 40128
rect 17868 39976 17920 39982
rect 17868 39918 17920 39924
rect 16500 39494 16712 39522
rect 16396 39432 16448 39438
rect 16396 39374 16448 39380
rect 16304 38956 16356 38962
rect 16304 38898 16356 38904
rect 15844 38344 15896 38350
rect 15844 38286 15896 38292
rect 16212 38344 16264 38350
rect 16212 38286 16264 38292
rect 15660 38208 15712 38214
rect 15660 38150 15712 38156
rect 15672 37874 15700 38150
rect 15568 37868 15620 37874
rect 15568 37810 15620 37816
rect 15660 37868 15712 37874
rect 15660 37810 15712 37816
rect 15476 37732 15528 37738
rect 15476 37674 15528 37680
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15108 35488 15160 35494
rect 15108 35430 15160 35436
rect 14924 34944 14976 34950
rect 14924 34886 14976 34892
rect 14740 34740 14792 34746
rect 14740 34682 14792 34688
rect 14936 34610 14964 34886
rect 15120 34610 15148 35430
rect 15384 34672 15436 34678
rect 15384 34614 15436 34620
rect 14188 34604 14240 34610
rect 14188 34546 14240 34552
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14924 34604 14976 34610
rect 14924 34546 14976 34552
rect 15108 34604 15160 34610
rect 15108 34546 15160 34552
rect 14200 33522 14228 34546
rect 14660 33998 14688 34546
rect 15396 34474 15424 34614
rect 15580 34610 15608 37810
rect 15568 34604 15620 34610
rect 15568 34546 15620 34552
rect 15384 34468 15436 34474
rect 15384 34410 15436 34416
rect 15292 34400 15344 34406
rect 15292 34342 15344 34348
rect 14372 33992 14424 33998
rect 14372 33934 14424 33940
rect 14648 33992 14700 33998
rect 14648 33934 14700 33940
rect 15016 33992 15068 33998
rect 15016 33934 15068 33940
rect 14188 33516 14240 33522
rect 14188 33458 14240 33464
rect 14096 33380 14148 33386
rect 14096 33322 14148 33328
rect 13912 33312 13964 33318
rect 13912 33254 13964 33260
rect 13820 32972 13872 32978
rect 13820 32914 13872 32920
rect 13832 32502 13860 32914
rect 13924 32910 13952 33254
rect 14108 32910 14136 33322
rect 13912 32904 13964 32910
rect 13912 32846 13964 32852
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 13820 32496 13872 32502
rect 13820 32438 13872 32444
rect 14200 32298 14228 33458
rect 14280 33448 14332 33454
rect 14280 33390 14332 33396
rect 14292 32910 14320 33390
rect 14280 32904 14332 32910
rect 14280 32846 14332 32852
rect 14384 32842 14412 33934
rect 14556 33856 14608 33862
rect 14556 33798 14608 33804
rect 14568 33590 14596 33798
rect 14556 33584 14608 33590
rect 14556 33526 14608 33532
rect 15028 33522 15056 33934
rect 15304 33930 15332 34342
rect 15292 33924 15344 33930
rect 15292 33866 15344 33872
rect 14464 33516 14516 33522
rect 14464 33458 14516 33464
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 14476 33114 14504 33458
rect 14464 33108 14516 33114
rect 14464 33050 14516 33056
rect 15028 32978 15056 33458
rect 15016 32972 15068 32978
rect 15016 32914 15068 32920
rect 14372 32836 14424 32842
rect 14372 32778 14424 32784
rect 15028 32434 15056 32914
rect 15016 32428 15068 32434
rect 15016 32370 15068 32376
rect 15292 32428 15344 32434
rect 15292 32370 15344 32376
rect 14188 32292 14240 32298
rect 14188 32234 14240 32240
rect 15304 32026 15332 32370
rect 15292 32020 15344 32026
rect 15292 31962 15344 31968
rect 15108 29844 15160 29850
rect 15108 29786 15160 29792
rect 13544 29232 13596 29238
rect 13544 29174 13596 29180
rect 15120 29170 15148 29786
rect 12992 29164 13044 29170
rect 12992 29106 13044 29112
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13820 29164 13872 29170
rect 13820 29106 13872 29112
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 15292 29164 15344 29170
rect 15292 29106 15344 29112
rect 13004 28762 13032 29106
rect 12992 28756 13044 28762
rect 12992 28698 13044 28704
rect 13004 27130 13032 28698
rect 13084 28620 13136 28626
rect 13084 28562 13136 28568
rect 13096 28218 13124 28562
rect 13648 28422 13676 29106
rect 13832 28490 13860 29106
rect 15200 29096 15252 29102
rect 15200 29038 15252 29044
rect 14372 29028 14424 29034
rect 14372 28970 14424 28976
rect 14740 29028 14792 29034
rect 14740 28970 14792 28976
rect 14096 28552 14148 28558
rect 14096 28494 14148 28500
rect 13820 28484 13872 28490
rect 13820 28426 13872 28432
rect 13636 28416 13688 28422
rect 13636 28358 13688 28364
rect 13084 28212 13136 28218
rect 13084 28154 13136 28160
rect 13096 27538 13124 28154
rect 13360 28008 13412 28014
rect 13360 27950 13412 27956
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 12992 27124 13044 27130
rect 12992 27066 13044 27072
rect 13096 26994 13124 27474
rect 13084 26988 13136 26994
rect 13084 26930 13136 26936
rect 13372 26042 13400 27950
rect 13648 26790 13676 28358
rect 13832 26994 13860 28426
rect 14004 27940 14056 27946
rect 14004 27882 14056 27888
rect 13912 27056 13964 27062
rect 13912 26998 13964 27004
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13832 26586 13860 26930
rect 13820 26580 13872 26586
rect 13820 26522 13872 26528
rect 13360 26036 13412 26042
rect 13360 25978 13412 25984
rect 13924 25838 13952 26998
rect 14016 26994 14044 27882
rect 14108 27538 14136 28494
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 14200 27674 14228 28086
rect 14188 27668 14240 27674
rect 14188 27610 14240 27616
rect 14096 27532 14148 27538
rect 14096 27474 14148 27480
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 14384 26926 14412 28970
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14660 27062 14688 28494
rect 14648 27056 14700 27062
rect 14648 26998 14700 27004
rect 14752 26994 14780 28970
rect 15212 27402 15240 29038
rect 15304 28762 15332 29106
rect 15292 28756 15344 28762
rect 15292 28698 15344 28704
rect 15396 28218 15424 34410
rect 15580 33658 15608 34546
rect 15856 34202 15884 38286
rect 16120 38276 16172 38282
rect 16120 38218 16172 38224
rect 16132 37942 16160 38218
rect 16120 37936 16172 37942
rect 16120 37878 16172 37884
rect 15936 37800 15988 37806
rect 15936 37742 15988 37748
rect 15948 37194 15976 37742
rect 15936 37188 15988 37194
rect 15936 37130 15988 37136
rect 15948 36786 15976 37130
rect 16212 36848 16264 36854
rect 16212 36790 16264 36796
rect 15936 36780 15988 36786
rect 15936 36722 15988 36728
rect 15948 36666 15976 36722
rect 15948 36638 16068 36666
rect 16040 36582 16068 36638
rect 16028 36576 16080 36582
rect 16028 36518 16080 36524
rect 16224 35834 16252 36790
rect 16212 35828 16264 35834
rect 16212 35770 16264 35776
rect 16224 34746 16252 35770
rect 16304 35692 16356 35698
rect 16304 35634 16356 35640
rect 16316 34950 16344 35634
rect 16408 35290 16436 39374
rect 16488 39364 16540 39370
rect 16488 39306 16540 39312
rect 16500 38706 16528 39306
rect 16500 38678 16620 38706
rect 16488 38412 16540 38418
rect 16488 38354 16540 38360
rect 16500 37466 16528 38354
rect 16592 38282 16620 38678
rect 16684 38332 16712 39494
rect 16856 39296 16908 39302
rect 16856 39238 16908 39244
rect 16868 38962 16896 39238
rect 17880 39098 17908 39918
rect 17868 39092 17920 39098
rect 17868 39034 17920 39040
rect 16856 38956 16908 38962
rect 16856 38898 16908 38904
rect 16868 38554 16896 38898
rect 18156 38894 18184 44678
rect 18432 44470 18460 44814
rect 18236 44464 18288 44470
rect 18236 44406 18288 44412
rect 18420 44464 18472 44470
rect 18420 44406 18472 44412
rect 18248 43314 18276 44406
rect 19352 43926 19380 44814
rect 19536 44266 19564 45426
rect 19996 45082 20024 45426
rect 19984 45076 20036 45082
rect 19984 45018 20036 45024
rect 20640 44402 20668 45494
rect 22112 45354 22140 46990
rect 22100 45348 22152 45354
rect 22100 45290 22152 45296
rect 20628 44396 20680 44402
rect 20628 44338 20680 44344
rect 19524 44260 19576 44266
rect 19524 44202 19576 44208
rect 20076 44192 20128 44198
rect 20076 44134 20128 44140
rect 19340 43920 19392 43926
rect 19340 43862 19392 43868
rect 19708 43784 19760 43790
rect 19708 43726 19760 43732
rect 19248 43648 19300 43654
rect 19248 43590 19300 43596
rect 18420 43444 18472 43450
rect 18420 43386 18472 43392
rect 18236 43308 18288 43314
rect 18236 43250 18288 43256
rect 18144 38888 18196 38894
rect 18144 38830 18196 38836
rect 18248 38758 18276 43250
rect 18432 42770 18460 43386
rect 19260 42770 19288 43590
rect 19340 43308 19392 43314
rect 19340 43250 19392 43256
rect 19352 42770 19380 43250
rect 19720 43110 19748 43726
rect 20088 43722 20116 44134
rect 20640 43994 20668 44338
rect 21180 44192 21232 44198
rect 21180 44134 21232 44140
rect 20260 43988 20312 43994
rect 20260 43930 20312 43936
rect 20628 43988 20680 43994
rect 20628 43930 20680 43936
rect 20076 43716 20128 43722
rect 20076 43658 20128 43664
rect 20272 43450 20300 43930
rect 20640 43790 20668 43930
rect 20628 43784 20680 43790
rect 20628 43726 20680 43732
rect 21192 43654 21220 44134
rect 21180 43648 21232 43654
rect 21180 43590 21232 43596
rect 20260 43444 20312 43450
rect 20260 43386 20312 43392
rect 19708 43104 19760 43110
rect 19708 43046 19760 43052
rect 18420 42764 18472 42770
rect 18420 42706 18472 42712
rect 19248 42764 19300 42770
rect 19248 42706 19300 42712
rect 19340 42764 19392 42770
rect 19340 42706 19392 42712
rect 19260 42650 19288 42706
rect 19432 42696 19484 42702
rect 19260 42622 19380 42650
rect 19432 42638 19484 42644
rect 18420 39840 18472 39846
rect 18420 39782 18472 39788
rect 18432 39438 18460 39782
rect 18420 39432 18472 39438
rect 18420 39374 18472 39380
rect 18696 39432 18748 39438
rect 18696 39374 18748 39380
rect 18708 39098 18736 39374
rect 19156 39296 19208 39302
rect 19156 39238 19208 39244
rect 18696 39092 18748 39098
rect 18696 39034 18748 39040
rect 19168 38962 19196 39238
rect 19156 38956 19208 38962
rect 19156 38898 19208 38904
rect 17592 38752 17644 38758
rect 17592 38694 17644 38700
rect 18236 38752 18288 38758
rect 18236 38694 18288 38700
rect 16856 38548 16908 38554
rect 16856 38490 16908 38496
rect 16868 38418 16896 38490
rect 17604 38418 17632 38694
rect 19352 38554 19380 42622
rect 19444 42362 19472 42638
rect 19432 42356 19484 42362
rect 19432 42298 19484 42304
rect 19720 42294 19748 43046
rect 19708 42288 19760 42294
rect 19708 42230 19760 42236
rect 21192 42022 21220 43590
rect 20168 42016 20220 42022
rect 20168 41958 20220 41964
rect 21180 42016 21232 42022
rect 21180 41958 21232 41964
rect 19524 39500 19576 39506
rect 19524 39442 19576 39448
rect 19536 38962 19564 39442
rect 19800 39024 19852 39030
rect 19800 38966 19852 38972
rect 19524 38956 19576 38962
rect 19524 38898 19576 38904
rect 19536 38842 19564 38898
rect 19444 38814 19564 38842
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 16856 38412 16908 38418
rect 16856 38354 16908 38360
rect 17592 38412 17644 38418
rect 17592 38354 17644 38360
rect 16764 38344 16816 38350
rect 16684 38304 16764 38332
rect 16764 38286 16816 38292
rect 16580 38276 16632 38282
rect 16580 38218 16632 38224
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16580 36916 16632 36922
rect 16580 36858 16632 36864
rect 16396 35284 16448 35290
rect 16396 35226 16448 35232
rect 16304 34944 16356 34950
rect 16304 34886 16356 34892
rect 16212 34740 16264 34746
rect 16212 34682 16264 34688
rect 16408 34678 16436 35226
rect 16592 35086 16620 36858
rect 16776 35834 16804 38286
rect 17316 37800 17368 37806
rect 17316 37742 17368 37748
rect 17328 36650 17356 37742
rect 17604 37330 17632 38354
rect 18604 38276 18656 38282
rect 18604 38218 18656 38224
rect 17776 38208 17828 38214
rect 17828 38168 17908 38196
rect 17776 38150 17828 38156
rect 17880 37806 17908 38168
rect 18616 38010 18644 38218
rect 19444 38010 19472 38814
rect 19524 38752 19576 38758
rect 19524 38694 19576 38700
rect 18604 38004 18656 38010
rect 18604 37946 18656 37952
rect 19432 38004 19484 38010
rect 19432 37946 19484 37952
rect 17868 37800 17920 37806
rect 17868 37742 17920 37748
rect 18420 37800 18472 37806
rect 18420 37742 18472 37748
rect 17684 37664 17736 37670
rect 17684 37606 17736 37612
rect 17592 37324 17644 37330
rect 17592 37266 17644 37272
rect 17696 37262 17724 37606
rect 17880 37466 17908 37742
rect 18432 37466 18460 37742
rect 17868 37460 17920 37466
rect 17868 37402 17920 37408
rect 18420 37460 18472 37466
rect 18420 37402 18472 37408
rect 17684 37256 17736 37262
rect 17684 37198 17736 37204
rect 17880 36922 17908 37402
rect 19536 37262 19564 38694
rect 19812 38350 19840 38966
rect 20180 38962 20208 41958
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 20168 38956 20220 38962
rect 20168 38898 20220 38904
rect 19996 38554 20024 38898
rect 23112 38752 23164 38758
rect 23112 38694 23164 38700
rect 19984 38548 20036 38554
rect 19984 38490 20036 38496
rect 19800 38344 19852 38350
rect 19800 38286 19852 38292
rect 19892 38208 19944 38214
rect 19892 38150 19944 38156
rect 19904 37806 19932 38150
rect 19892 37800 19944 37806
rect 19892 37742 19944 37748
rect 19904 37330 19932 37742
rect 19892 37324 19944 37330
rect 19892 37266 19944 37272
rect 19524 37256 19576 37262
rect 19524 37198 19576 37204
rect 17868 36916 17920 36922
rect 17868 36858 17920 36864
rect 17316 36644 17368 36650
rect 17316 36586 17368 36592
rect 23124 35894 23152 38694
rect 23124 35866 23244 35894
rect 16764 35828 16816 35834
rect 16764 35770 16816 35776
rect 16776 35222 16804 35770
rect 16764 35216 16816 35222
rect 16764 35158 16816 35164
rect 17592 35216 17644 35222
rect 17592 35158 17644 35164
rect 16580 35080 16632 35086
rect 16580 35022 16632 35028
rect 16396 34672 16448 34678
rect 16396 34614 16448 34620
rect 16592 34202 16620 35022
rect 15844 34196 15896 34202
rect 15844 34138 15896 34144
rect 16580 34196 16632 34202
rect 16580 34138 16632 34144
rect 15568 33652 15620 33658
rect 15568 33594 15620 33600
rect 16776 33114 16804 35158
rect 17604 34066 17632 35158
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 17868 34400 17920 34406
rect 17868 34342 17920 34348
rect 18788 34400 18840 34406
rect 18788 34342 18840 34348
rect 17592 34060 17644 34066
rect 17592 34002 17644 34008
rect 17684 33992 17736 33998
rect 17880 33980 17908 34342
rect 18800 34202 18828 34342
rect 18788 34196 18840 34202
rect 18788 34138 18840 34144
rect 17736 33952 17908 33980
rect 17684 33934 17736 33940
rect 17500 33924 17552 33930
rect 17500 33866 17552 33872
rect 17512 33114 17540 33866
rect 17880 33590 17908 33952
rect 19156 33992 19208 33998
rect 19156 33934 19208 33940
rect 18052 33856 18104 33862
rect 18052 33798 18104 33804
rect 17868 33584 17920 33590
rect 17868 33526 17920 33532
rect 18064 33522 18092 33798
rect 19168 33658 19196 33934
rect 19340 33856 19392 33862
rect 19340 33798 19392 33804
rect 19156 33652 19208 33658
rect 19156 33594 19208 33600
rect 17592 33516 17644 33522
rect 17592 33458 17644 33464
rect 18052 33516 18104 33522
rect 18052 33458 18104 33464
rect 16764 33108 16816 33114
rect 16764 33050 16816 33056
rect 17500 33108 17552 33114
rect 17500 33050 17552 33056
rect 16488 33040 16540 33046
rect 16488 32982 16540 32988
rect 15752 32768 15804 32774
rect 15752 32710 15804 32716
rect 15764 32570 15792 32710
rect 15752 32564 15804 32570
rect 15752 32506 15804 32512
rect 16396 32564 16448 32570
rect 16396 32506 16448 32512
rect 16408 31890 16436 32506
rect 16396 31884 16448 31890
rect 16396 31826 16448 31832
rect 16408 29170 16436 31826
rect 16500 31822 16528 32982
rect 16776 32842 16804 33050
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 17040 32496 17092 32502
rect 17040 32438 17092 32444
rect 17052 32026 17080 32438
rect 17040 32020 17092 32026
rect 17040 31962 17092 31968
rect 16488 31816 16540 31822
rect 16488 31758 16540 31764
rect 16396 29164 16448 29170
rect 16396 29106 16448 29112
rect 16764 29164 16816 29170
rect 16948 29164 17000 29170
rect 16816 29124 16896 29152
rect 16764 29106 16816 29112
rect 16764 29028 16816 29034
rect 16764 28970 16816 28976
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 15384 28212 15436 28218
rect 15384 28154 15436 28160
rect 16592 27606 16620 28494
rect 16684 28082 16712 28494
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16580 27600 16632 27606
rect 16580 27542 16632 27548
rect 16684 27402 16712 28018
rect 16776 27538 16804 28970
rect 16868 28762 16896 29124
rect 16948 29106 17000 29112
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 16960 28218 16988 29106
rect 17052 28966 17080 31962
rect 17316 30116 17368 30122
rect 17316 30058 17368 30064
rect 17328 29850 17356 30058
rect 17500 30048 17552 30054
rect 17500 29990 17552 29996
rect 17316 29844 17368 29850
rect 17316 29786 17368 29792
rect 17512 29646 17540 29990
rect 17604 29714 17632 33458
rect 19352 33114 19380 33798
rect 19444 33658 19472 34478
rect 22192 33992 22244 33998
rect 22192 33934 22244 33940
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 21548 33856 21600 33862
rect 21548 33798 21600 33804
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 19996 33522 20024 33798
rect 21560 33522 21588 33798
rect 19984 33516 20036 33522
rect 19984 33458 20036 33464
rect 21548 33516 21600 33522
rect 21548 33458 21600 33464
rect 19708 33448 19760 33454
rect 19708 33390 19760 33396
rect 19340 33108 19392 33114
rect 19340 33050 19392 33056
rect 19720 33046 19748 33390
rect 19708 33040 19760 33046
rect 19628 32988 19708 32994
rect 19628 32982 19760 32988
rect 18880 32972 18932 32978
rect 18880 32914 18932 32920
rect 19628 32966 19748 32982
rect 17684 32904 17736 32910
rect 17684 32846 17736 32852
rect 17696 32570 17724 32846
rect 17776 32836 17828 32842
rect 17776 32778 17828 32784
rect 17684 32564 17736 32570
rect 17684 32506 17736 32512
rect 17684 30660 17736 30666
rect 17684 30602 17736 30608
rect 17696 30258 17724 30602
rect 17788 30598 17816 32778
rect 18604 32768 18656 32774
rect 18604 32710 18656 32716
rect 18616 32026 18644 32710
rect 18892 32434 18920 32914
rect 19628 32570 19656 32966
rect 19996 32910 20024 33458
rect 22204 33114 22232 33934
rect 22192 33108 22244 33114
rect 22192 33050 22244 33056
rect 21180 32972 21232 32978
rect 21180 32914 21232 32920
rect 19708 32904 19760 32910
rect 19708 32846 19760 32852
rect 19984 32904 20036 32910
rect 19984 32846 20036 32852
rect 19616 32564 19668 32570
rect 19616 32506 19668 32512
rect 18880 32428 18932 32434
rect 18880 32370 18932 32376
rect 18788 32224 18840 32230
rect 18788 32166 18840 32172
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 18800 31822 18828 32166
rect 18892 31822 18920 32370
rect 19432 32292 19484 32298
rect 19432 32234 19484 32240
rect 19248 31884 19300 31890
rect 19248 31826 19300 31832
rect 18788 31816 18840 31822
rect 18788 31758 18840 31764
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18604 31748 18656 31754
rect 18604 31690 18656 31696
rect 18616 30938 18644 31690
rect 18604 30932 18656 30938
rect 18604 30874 18656 30880
rect 17776 30592 17828 30598
rect 17776 30534 17828 30540
rect 17684 30252 17736 30258
rect 17684 30194 17736 30200
rect 17592 29708 17644 29714
rect 17592 29650 17644 29656
rect 17500 29640 17552 29646
rect 17500 29582 17552 29588
rect 17040 28960 17092 28966
rect 17040 28902 17092 28908
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 17052 27538 17080 28902
rect 17500 28756 17552 28762
rect 17500 28698 17552 28704
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 16764 27532 16816 27538
rect 16764 27474 16816 27480
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 16856 27464 16908 27470
rect 16856 27406 16908 27412
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 16672 27396 16724 27402
rect 16672 27338 16724 27344
rect 16684 27130 16712 27338
rect 16764 27328 16816 27334
rect 16764 27270 16816 27276
rect 16672 27124 16724 27130
rect 16672 27066 16724 27072
rect 16776 26994 16804 27270
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16868 26926 16896 27406
rect 14372 26920 14424 26926
rect 14372 26862 14424 26868
rect 16856 26920 16908 26926
rect 16856 26862 16908 26868
rect 17052 26858 17080 27474
rect 17144 27470 17172 28494
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 17224 27940 17276 27946
rect 17224 27882 17276 27888
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17040 26852 17092 26858
rect 17040 26794 17092 26800
rect 17144 26382 17172 27270
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 17040 26308 17092 26314
rect 17040 26250 17092 26256
rect 13912 25832 13964 25838
rect 13912 25774 13964 25780
rect 13924 24682 13952 25774
rect 13912 24676 13964 24682
rect 13912 24618 13964 24624
rect 17052 24274 17080 26250
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16316 23798 16344 24006
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 14464 23724 14516 23730
rect 14464 23666 14516 23672
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 13544 23588 13596 23594
rect 13544 23530 13596 23536
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 13280 23118 13308 23462
rect 13556 23254 13584 23530
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13544 23248 13596 23254
rect 13544 23190 13596 23196
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13556 21962 13584 23190
rect 13648 22710 13676 23462
rect 13728 23180 13780 23186
rect 13728 23122 13780 23128
rect 14004 23180 14056 23186
rect 14004 23122 14056 23128
rect 13636 22704 13688 22710
rect 13636 22646 13688 22652
rect 13740 21962 13768 23122
rect 14016 22574 14044 23122
rect 14292 22778 14320 23598
rect 14476 23118 14504 23666
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15672 23118 15700 23462
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 14016 22030 14044 22510
rect 14660 22234 14688 23054
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13728 21956 13780 21962
rect 13728 21898 13780 21904
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9036 18896 9088 18902
rect 9036 18838 9088 18844
rect 9048 18766 9076 18838
rect 9232 18766 9260 19110
rect 9312 18896 9364 18902
rect 9312 18838 9364 18844
rect 7564 18760 7616 18766
rect 6920 18692 6972 18698
rect 7116 18686 7236 18714
rect 7564 18702 7616 18708
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 6920 18634 6972 18640
rect 6644 18624 6696 18630
rect 6644 18566 6696 18572
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5920 17202 5948 17478
rect 6104 17338 6132 17546
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6656 17202 6684 18566
rect 6748 18290 6776 18566
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6932 17338 6960 18634
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18426 7144 18566
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4724 16794 4752 16934
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 5644 16590 5672 17070
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 7024 16454 7052 18226
rect 7116 16658 7144 18362
rect 7208 17882 7236 18686
rect 7576 18086 7604 18702
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 7852 18426 7880 18634
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7208 16590 7236 17818
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7300 16590 7328 17274
rect 7852 16658 7880 18362
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 8220 17882 8248 18158
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 9324 17678 9352 18838
rect 9416 18630 9444 19314
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 9968 18766 9996 18906
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9416 18426 9444 18566
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9416 17746 9444 18362
rect 9600 18358 9628 18702
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 8036 17270 8064 17614
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 9416 17202 9444 17682
rect 9508 17678 9536 17818
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9508 17542 9536 17614
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9600 17338 9628 18294
rect 10060 18154 10088 19246
rect 10520 18970 10548 19246
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 10152 17270 10180 18022
rect 10612 17882 10640 19314
rect 10888 18834 10916 19382
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10704 18222 10732 18566
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10140 17264 10192 17270
rect 10140 17206 10192 17212
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 8220 16794 8248 17138
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 10980 16726 11008 18566
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 9784 15026 9812 15438
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10980 15162 11008 15370
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 7116 13870 7144 14418
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 6932 12918 6960 13670
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 7024 12986 7052 13194
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5460 11218 5488 12174
rect 5552 11762 5580 12786
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 12170 5764 12582
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 6104 11898 6132 12718
rect 7116 12434 7144 13806
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7300 12850 7328 13262
rect 7392 12918 7420 14282
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7576 12918 7604 14214
rect 7944 14074 7972 14350
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8128 13530 8156 13806
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7564 12912 7616 12918
rect 7564 12854 7616 12860
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7024 12406 7144 12434
rect 7024 12102 7052 12406
rect 7300 12238 7328 12786
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5736 11150 5764 11494
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5920 2650 5948 11698
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 11354 6868 11630
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 7024 11286 7052 12038
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7392 11150 7420 12854
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7944 11354 7972 12106
rect 8312 11898 8340 14282
rect 8404 12986 8432 14350
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8312 11762 8340 11834
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8312 11642 8340 11698
rect 8496 11694 8524 14554
rect 9692 14278 9720 14894
rect 9784 14618 9812 14962
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 13410 9720 14214
rect 9784 13530 9812 14554
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9600 13382 9720 13410
rect 10152 13394 10180 13874
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10140 13388 10192 13394
rect 9600 13326 9628 13382
rect 10140 13330 10192 13336
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9140 12986 9168 13262
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 8484 11688 8536 11694
rect 8312 11614 8432 11642
rect 8484 11630 8536 11636
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 8312 11218 8340 11494
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8404 11150 8432 11614
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8496 11082 8524 11630
rect 9416 11150 9444 12378
rect 9600 11150 9628 13262
rect 9692 11354 9720 13262
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 9968 12918 9996 13126
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 10152 12434 10180 13126
rect 10244 12850 10272 13670
rect 10336 13530 10364 13806
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10612 13394 10640 13874
rect 10980 13870 11008 15098
rect 11348 14618 11376 18226
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11624 15026 11652 17818
rect 11808 17678 11836 18022
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11716 16658 11744 17274
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11716 15502 11744 16594
rect 11808 16114 11836 17614
rect 11900 16726 11928 17614
rect 12176 17338 12204 18158
rect 12268 17678 12296 20402
rect 13464 19514 13492 21490
rect 13740 21146 13768 21898
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 14016 20398 14044 21966
rect 15764 21010 15792 23666
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16776 23322 16804 23598
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 17052 23254 17080 24210
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 17236 21962 17264 27882
rect 17420 27130 17448 27950
rect 17512 27606 17540 28698
rect 17604 27674 17632 29650
rect 17696 28694 17724 30194
rect 17788 30122 17816 30534
rect 18616 30326 18644 30874
rect 18604 30320 18656 30326
rect 18604 30262 18656 30268
rect 17776 30116 17828 30122
rect 17776 30058 17828 30064
rect 18604 30048 18656 30054
rect 18604 29990 18656 29996
rect 18616 29714 18644 29990
rect 18800 29850 18828 31758
rect 19260 30734 19288 31826
rect 19444 31822 19472 32234
rect 19720 31890 19748 32846
rect 19996 32434 20024 32846
rect 20168 32768 20220 32774
rect 20168 32710 20220 32716
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19708 31884 19760 31890
rect 19708 31826 19760 31832
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19616 31816 19668 31822
rect 19616 31758 19668 31764
rect 19628 30802 19656 31758
rect 19616 30796 19668 30802
rect 19616 30738 19668 30744
rect 19248 30728 19300 30734
rect 19248 30670 19300 30676
rect 19628 30258 19656 30738
rect 19616 30252 19668 30258
rect 19616 30194 19668 30200
rect 19340 30184 19392 30190
rect 19340 30126 19392 30132
rect 19352 29850 19380 30126
rect 18788 29844 18840 29850
rect 18788 29786 18840 29792
rect 19340 29844 19392 29850
rect 19340 29786 19392 29792
rect 18604 29708 18656 29714
rect 18604 29650 18656 29656
rect 18144 29232 18196 29238
rect 18144 29174 18196 29180
rect 17960 29096 18012 29102
rect 17960 29038 18012 29044
rect 17684 28688 17736 28694
rect 17684 28630 17736 28636
rect 17776 28552 17828 28558
rect 17776 28494 17828 28500
rect 17684 28484 17736 28490
rect 17684 28426 17736 28432
rect 17696 28082 17724 28426
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17696 27674 17724 28018
rect 17592 27668 17644 27674
rect 17592 27610 17644 27616
rect 17684 27668 17736 27674
rect 17684 27610 17736 27616
rect 17500 27600 17552 27606
rect 17500 27542 17552 27548
rect 17788 27334 17816 28494
rect 17972 28082 18000 29038
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 18156 27470 18184 29174
rect 18800 29170 18828 29786
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 18788 29164 18840 29170
rect 18788 29106 18840 29112
rect 19444 29102 19472 29446
rect 19628 29306 19656 30194
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19616 29300 19668 29306
rect 19616 29242 19668 29248
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 19444 28422 19472 29038
rect 19904 29034 19932 29650
rect 19892 29028 19944 29034
rect 19892 28970 19944 28976
rect 19524 28960 19576 28966
rect 19524 28902 19576 28908
rect 19536 28558 19564 28902
rect 19904 28558 19932 28970
rect 19524 28552 19576 28558
rect 19524 28494 19576 28500
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 17868 27396 17920 27402
rect 17868 27338 17920 27344
rect 17776 27328 17828 27334
rect 17776 27270 17828 27276
rect 17408 27124 17460 27130
rect 17408 27066 17460 27072
rect 17684 26920 17736 26926
rect 17684 26862 17736 26868
rect 17696 26586 17724 26862
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 17880 26314 17908 27338
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 17972 26586 18000 26930
rect 17960 26580 18012 26586
rect 17960 26522 18012 26528
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17316 24064 17368 24070
rect 17316 24006 17368 24012
rect 17328 23798 17356 24006
rect 17512 23866 17540 24142
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17316 23792 17368 23798
rect 17316 23734 17368 23740
rect 17604 23730 17632 24142
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17972 23050 18000 24550
rect 18064 24206 18092 24822
rect 18156 24206 18184 26318
rect 18616 26042 18644 26930
rect 19156 26444 19208 26450
rect 19156 26386 19208 26392
rect 18604 26036 18656 26042
rect 18604 25978 18656 25984
rect 19168 25906 19196 26386
rect 19444 26382 19472 28358
rect 19892 26784 19944 26790
rect 19892 26726 19944 26732
rect 19904 26382 19932 26726
rect 20180 26450 20208 32710
rect 21192 32026 21220 32914
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 21928 32570 21956 32846
rect 21916 32564 21968 32570
rect 21916 32506 21968 32512
rect 21928 32450 21956 32506
rect 21928 32422 22140 32450
rect 22388 32434 22416 32846
rect 21916 32360 21968 32366
rect 21916 32302 21968 32308
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 21180 32020 21232 32026
rect 21180 31962 21232 31968
rect 21100 31822 21128 31962
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 21456 31816 21508 31822
rect 21456 31758 21508 31764
rect 20812 31748 20864 31754
rect 20812 31690 20864 31696
rect 21180 31748 21232 31754
rect 21180 31690 21232 31696
rect 20824 31414 20852 31690
rect 20812 31408 20864 31414
rect 20812 31350 20864 31356
rect 21192 31346 21220 31690
rect 21180 31340 21232 31346
rect 21180 31282 21232 31288
rect 21468 31278 21496 31758
rect 21928 31414 21956 32302
rect 22112 31822 22140 32422
rect 22376 32428 22428 32434
rect 22376 32370 22428 32376
rect 22192 32224 22244 32230
rect 22192 32166 22244 32172
rect 22204 31890 22232 32166
rect 22192 31884 22244 31890
rect 22192 31826 22244 31832
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 21916 31408 21968 31414
rect 21916 31350 21968 31356
rect 21456 31272 21508 31278
rect 21456 31214 21508 31220
rect 21548 31204 21600 31210
rect 21548 31146 21600 31152
rect 20628 30116 20680 30122
rect 20628 30058 20680 30064
rect 20640 28014 20668 30058
rect 21560 28626 21588 31146
rect 21928 29714 21956 31350
rect 22020 31278 22048 31758
rect 22100 31680 22152 31686
rect 22100 31622 22152 31628
rect 22112 31414 22140 31622
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22008 31272 22060 31278
rect 22008 31214 22060 31220
rect 21916 29708 21968 29714
rect 21916 29650 21968 29656
rect 21928 29238 21956 29650
rect 21916 29232 21968 29238
rect 21916 29174 21968 29180
rect 21548 28620 21600 28626
rect 21548 28562 21600 28568
rect 20904 28416 20956 28422
rect 20904 28358 20956 28364
rect 21548 28416 21600 28422
rect 21548 28358 21600 28364
rect 20916 28082 20944 28358
rect 20904 28076 20956 28082
rect 20904 28018 20956 28024
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 21560 27878 21588 28358
rect 22112 28218 22140 31350
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 20904 27872 20956 27878
rect 20904 27814 20956 27820
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 22008 27872 22060 27878
rect 22008 27814 22060 27820
rect 20916 27402 20944 27814
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 20904 27396 20956 27402
rect 20904 27338 20956 27344
rect 20260 27056 20312 27062
rect 20260 26998 20312 27004
rect 20272 26450 20300 26998
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20640 26586 20668 26930
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20168 26444 20220 26450
rect 20168 26386 20220 26392
rect 20260 26444 20312 26450
rect 20260 26386 20312 26392
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19892 26376 19944 26382
rect 19892 26318 19944 26324
rect 19444 25906 19472 26318
rect 20180 25974 20208 26386
rect 20168 25968 20220 25974
rect 20168 25910 20220 25916
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18248 24274 18276 24754
rect 18512 24676 18564 24682
rect 18512 24618 18564 24624
rect 18236 24268 18288 24274
rect 18236 24210 18288 24216
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 17960 23044 18012 23050
rect 17960 22986 18012 22992
rect 17972 22710 18000 22986
rect 18064 22982 18092 24142
rect 18156 23866 18184 24142
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18156 23118 18184 23802
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 18420 22976 18472 22982
rect 18420 22918 18472 22924
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 18432 22642 18460 22918
rect 18524 22642 18552 24618
rect 18616 23526 18644 25774
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19524 25152 19576 25158
rect 19524 25094 19576 25100
rect 19536 24818 19564 25094
rect 19524 24812 19576 24818
rect 19524 24754 19576 24760
rect 19812 24614 19840 25230
rect 20076 24744 20128 24750
rect 20076 24686 20128 24692
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19800 24608 19852 24614
rect 19800 24550 19852 24556
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18616 22642 18644 23462
rect 18696 23112 18748 23118
rect 18696 23054 18748 23060
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18708 22234 18736 23054
rect 19352 22778 19380 24142
rect 19444 23050 19472 24550
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19536 23798 19564 24006
rect 19524 23792 19576 23798
rect 19524 23734 19576 23740
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19812 22778 19840 24550
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 20088 22642 20116 24686
rect 20272 24206 20300 26386
rect 21180 26308 21232 26314
rect 21180 26250 21232 26256
rect 21192 26042 21220 26250
rect 20996 26036 21048 26042
rect 20996 25978 21048 25984
rect 21180 26036 21232 26042
rect 21180 25978 21232 25984
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20260 24200 20312 24206
rect 20260 24142 20312 24148
rect 20272 23866 20300 24142
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20548 23118 20576 25230
rect 20904 25220 20956 25226
rect 20904 25162 20956 25168
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20732 24682 20760 25094
rect 20812 24744 20864 24750
rect 20916 24698 20944 25162
rect 21008 24750 21036 25978
rect 21180 25492 21232 25498
rect 21180 25434 21232 25440
rect 21192 24886 21220 25434
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 21180 24880 21232 24886
rect 21180 24822 21232 24828
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 20864 24692 20944 24698
rect 20812 24686 20944 24692
rect 20996 24744 21048 24750
rect 20996 24686 21048 24692
rect 20720 24676 20772 24682
rect 20824 24670 20944 24686
rect 20720 24618 20772 24624
rect 20628 24608 20680 24614
rect 20628 24550 20680 24556
rect 20640 24274 20668 24550
rect 20916 24410 20944 24670
rect 20904 24404 20956 24410
rect 20904 24346 20956 24352
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 21008 23322 21036 24686
rect 21100 23322 21128 24754
rect 21284 24682 21312 25094
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21284 24138 21312 24618
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21180 24064 21232 24070
rect 21180 24006 21232 24012
rect 21192 23730 21220 24006
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 21284 23118 21312 24074
rect 21468 23730 21496 27406
rect 22020 26994 22048 27814
rect 22204 27674 22232 28018
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 22388 27130 22416 32370
rect 23112 32224 23164 32230
rect 23112 32166 23164 32172
rect 22744 31816 22796 31822
rect 22744 31758 22796 31764
rect 22756 31482 22784 31758
rect 22744 31476 22796 31482
rect 22744 31418 22796 31424
rect 23124 28082 23152 32166
rect 23216 28558 23244 35866
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 24492 33856 24544 33862
rect 24492 33798 24544 33804
rect 24504 33590 24532 33798
rect 24492 33584 24544 33590
rect 24492 33526 24544 33532
rect 23756 33516 23808 33522
rect 23756 33458 23808 33464
rect 23572 33380 23624 33386
rect 23572 33322 23624 33328
rect 23296 33312 23348 33318
rect 23296 33254 23348 33260
rect 23308 32978 23336 33254
rect 23296 32972 23348 32978
rect 23296 32914 23348 32920
rect 23388 32972 23440 32978
rect 23388 32914 23440 32920
rect 23308 32434 23336 32914
rect 23400 32502 23428 32914
rect 23388 32496 23440 32502
rect 23388 32438 23440 32444
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 23584 32366 23612 33322
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23676 32910 23704 33254
rect 23768 33114 23796 33458
rect 23756 33108 23808 33114
rect 23756 33050 23808 33056
rect 23848 33040 23900 33046
rect 23848 32982 23900 32988
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23664 32768 23716 32774
rect 23664 32710 23716 32716
rect 23676 32434 23704 32710
rect 23860 32570 23888 32982
rect 24676 32768 24728 32774
rect 24676 32710 24728 32716
rect 23848 32564 23900 32570
rect 23848 32506 23900 32512
rect 23664 32428 23716 32434
rect 23664 32370 23716 32376
rect 23572 32360 23624 32366
rect 23572 32302 23624 32308
rect 23584 31822 23612 32302
rect 23860 32298 23888 32506
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 23848 32292 23900 32298
rect 23848 32234 23900 32240
rect 23756 32020 23808 32026
rect 23756 31962 23808 31968
rect 23572 31816 23624 31822
rect 23572 31758 23624 31764
rect 23768 30258 23796 31962
rect 24228 30326 24256 32370
rect 24688 32366 24716 32710
rect 24676 32360 24728 32366
rect 24676 32302 24728 32308
rect 25056 32230 25084 33934
rect 25320 33312 25372 33318
rect 25320 33254 25372 33260
rect 25688 33312 25740 33318
rect 25688 33254 25740 33260
rect 25136 32904 25188 32910
rect 25136 32846 25188 32852
rect 25148 32570 25176 32846
rect 25136 32564 25188 32570
rect 25136 32506 25188 32512
rect 25044 32224 25096 32230
rect 25044 32166 25096 32172
rect 25136 32224 25188 32230
rect 25136 32166 25188 32172
rect 24584 31816 24636 31822
rect 24584 31758 24636 31764
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 23756 30252 23808 30258
rect 23756 30194 23808 30200
rect 23848 30252 23900 30258
rect 23848 30194 23900 30200
rect 24124 30252 24176 30258
rect 24124 30194 24176 30200
rect 23768 29220 23796 30194
rect 23676 29192 23796 29220
rect 23676 29102 23704 29192
rect 23664 29096 23716 29102
rect 23664 29038 23716 29044
rect 23860 29034 23888 30194
rect 24136 29510 24164 30194
rect 24596 29850 24624 31758
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24124 29504 24176 29510
rect 24124 29446 24176 29452
rect 24136 29238 24164 29446
rect 24124 29232 24176 29238
rect 24124 29174 24176 29180
rect 23848 29028 23900 29034
rect 23848 28970 23900 28976
rect 24032 28960 24084 28966
rect 24032 28902 24084 28908
rect 23848 28620 23900 28626
rect 23848 28562 23900 28568
rect 23204 28552 23256 28558
rect 23204 28494 23256 28500
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23480 28416 23532 28422
rect 23480 28358 23532 28364
rect 23492 28082 23520 28358
rect 23112 28076 23164 28082
rect 23112 28018 23164 28024
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23480 27872 23532 27878
rect 23480 27814 23532 27820
rect 23492 27470 23520 27814
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 22376 27124 22428 27130
rect 22376 27066 22428 27072
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 22020 26382 22048 26930
rect 22284 26920 22336 26926
rect 22284 26862 22336 26868
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 22296 26314 22324 26862
rect 22388 26382 22416 27066
rect 23020 26988 23072 26994
rect 23020 26930 23072 26936
rect 23032 26586 23060 26930
rect 23020 26580 23072 26586
rect 23020 26522 23072 26528
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22284 26308 22336 26314
rect 22284 26250 22336 26256
rect 22836 26308 22888 26314
rect 22836 26250 22888 26256
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21468 23186 21496 23666
rect 21928 23662 21956 24550
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 21732 23520 21784 23526
rect 21732 23462 21784 23468
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 20548 22506 20576 23054
rect 21468 22642 21496 23122
rect 21744 23118 21772 23462
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 20536 22500 20588 22506
rect 20536 22442 20588 22448
rect 18696 22228 18748 22234
rect 18696 22170 18748 22176
rect 22112 22098 22140 24754
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22664 24274 22692 24550
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22652 24064 22704 24070
rect 22652 24006 22704 24012
rect 22664 22710 22692 24006
rect 22848 23662 22876 26250
rect 23388 24880 23440 24886
rect 23388 24822 23440 24828
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23124 24070 23152 24550
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22848 23322 22876 23598
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22652 22704 22704 22710
rect 22652 22646 22704 22652
rect 22100 22092 22152 22098
rect 22100 22034 22152 22040
rect 23124 22030 23152 24006
rect 23400 23322 23428 24822
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23584 24274 23612 24550
rect 23572 24268 23624 24274
rect 23572 24210 23624 24216
rect 23584 23866 23612 24210
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23388 23044 23440 23050
rect 23388 22986 23440 22992
rect 23400 22574 23428 22986
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23400 22030 23428 22510
rect 23676 22094 23704 28494
rect 23860 28014 23888 28562
rect 24044 28218 24072 28902
rect 24492 28552 24544 28558
rect 24492 28494 24544 28500
rect 24504 28218 24532 28494
rect 24596 28490 24624 29786
rect 24952 29572 25004 29578
rect 24952 29514 25004 29520
rect 24964 29306 24992 29514
rect 24952 29300 25004 29306
rect 24952 29242 25004 29248
rect 24860 28620 24912 28626
rect 24860 28562 24912 28568
rect 24584 28484 24636 28490
rect 24584 28426 24636 28432
rect 24596 28218 24624 28426
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 24492 28212 24544 28218
rect 24492 28154 24544 28160
rect 24584 28212 24636 28218
rect 24584 28154 24636 28160
rect 24032 28076 24084 28082
rect 24032 28018 24084 28024
rect 23848 28008 23900 28014
rect 23848 27950 23900 27956
rect 24044 27130 24072 28018
rect 24032 27124 24084 27130
rect 24032 27066 24084 27072
rect 24044 26994 24072 27066
rect 23940 26988 23992 26994
rect 23940 26930 23992 26936
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23768 24206 23796 24754
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23952 23186 23980 26930
rect 24872 26790 24900 28562
rect 24964 28082 24992 29242
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 24964 27674 24992 28018
rect 24952 27668 25004 27674
rect 24952 27610 25004 27616
rect 25148 27130 25176 32166
rect 25332 29170 25360 33254
rect 25700 32434 25728 33254
rect 25780 32904 25832 32910
rect 25780 32846 25832 32852
rect 25688 32428 25740 32434
rect 25688 32370 25740 32376
rect 25792 32230 25820 32846
rect 27068 32428 27120 32434
rect 27068 32370 27120 32376
rect 25780 32224 25832 32230
rect 25780 32166 25832 32172
rect 27080 29306 27108 32370
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28276 32065 28304 32302
rect 28262 32056 28318 32065
rect 28262 31991 28318 32000
rect 28448 31816 28500 31822
rect 28448 31758 28500 31764
rect 28460 31385 28488 31758
rect 28446 31376 28502 31385
rect 28446 31311 28502 31320
rect 27068 29300 27120 29306
rect 27068 29242 27120 29248
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 26056 29164 26108 29170
rect 26056 29106 26108 29112
rect 26068 28762 26096 29106
rect 26056 28756 26108 28762
rect 26056 28698 26108 28704
rect 28448 27464 28500 27470
rect 28448 27406 28500 27412
rect 28460 27305 28488 27406
rect 28446 27296 28502 27305
rect 28446 27231 28502 27240
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 25228 26988 25280 26994
rect 25228 26930 25280 26936
rect 25240 26858 25268 26930
rect 25228 26852 25280 26858
rect 25228 26794 25280 26800
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24952 26784 25004 26790
rect 24952 26726 25004 26732
rect 24964 25786 24992 26726
rect 24872 25758 24992 25786
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 23940 23180 23992 23186
rect 23940 23122 23992 23128
rect 23952 22778 23980 23122
rect 24136 22778 24164 24686
rect 24492 24608 24544 24614
rect 24492 24550 24544 24556
rect 24504 24206 24532 24550
rect 24676 24336 24728 24342
rect 24676 24278 24728 24284
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24308 24132 24360 24138
rect 24308 24074 24360 24080
rect 23940 22772 23992 22778
rect 23940 22714 23992 22720
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 23676 22066 23796 22094
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 15752 21004 15804 21010
rect 15752 20946 15804 20952
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 15028 20534 15056 20742
rect 15016 20528 15068 20534
rect 15016 20470 15068 20476
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14568 19922 14596 20334
rect 15580 20262 15608 20878
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 15028 19514 15056 19722
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12452 17202 12480 17750
rect 15212 17678 15240 20198
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15580 19378 15608 19926
rect 15764 19786 15792 20946
rect 16396 20868 16448 20874
rect 16396 20810 16448 20816
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15764 19446 15792 19722
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 16040 19378 16068 19858
rect 16408 19854 16436 20810
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15660 19304 15712 19310
rect 15660 19246 15712 19252
rect 15672 18290 15700 19246
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18834 15884 19110
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15396 17678 15424 18158
rect 16040 18086 16068 19314
rect 16316 19310 16344 19654
rect 16408 19446 16436 19790
rect 16396 19440 16448 19446
rect 16396 19382 16448 19388
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16224 18358 16252 19246
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16316 18222 16344 19246
rect 16408 18358 16436 19382
rect 16500 19378 16528 19790
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16684 18358 16712 19178
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16776 18086 16804 18158
rect 16868 18154 16896 21830
rect 19892 20528 19944 20534
rect 19892 20470 19944 20476
rect 21824 20528 21876 20534
rect 21824 20470 21876 20476
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18156 19854 18184 19994
rect 19904 19922 19932 20470
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18156 19718 18184 19790
rect 18340 19718 18368 19790
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 17420 18698 17448 19654
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18156 18766 18184 19246
rect 18984 18970 19012 19790
rect 19996 19786 20024 20198
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 18970 19472 19654
rect 20272 19378 20300 20402
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 21100 20058 21128 20334
rect 21192 20262 21220 20402
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17882 16804 18022
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 17328 17746 17356 18566
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 11888 16720 11940 16726
rect 11888 16662 11940 16668
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11900 16046 11928 16526
rect 12268 16522 12296 17138
rect 12452 16590 12480 17138
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11900 15026 11928 15982
rect 12268 15570 12296 16458
rect 12452 15706 12480 16526
rect 12544 16250 12572 16594
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 13188 16114 13216 16390
rect 13280 16114 13308 16934
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13648 15706 13676 16186
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 13648 15502 13676 15642
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14618 11928 14962
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11348 14414 11376 14554
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10152 12406 10272 12434
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9968 11762 9996 12174
rect 10244 12170 10272 12406
rect 10612 12238 10640 13330
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12986 10916 13194
rect 11348 12986 11376 13262
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11348 12442 11376 12922
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11624 12442 11652 12718
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9588 11144 9640 11150
rect 9640 11092 9720 11098
rect 9588 11086 9720 11092
rect 8484 11076 8536 11082
rect 9600 11070 9720 11086
rect 8484 11018 8536 11024
rect 9692 10674 9720 11070
rect 9876 10810 9904 11698
rect 10060 11218 10088 12038
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 10612 10674 10640 11494
rect 10704 11354 10732 12106
rect 11348 11762 11376 12378
rect 12452 12238 12480 13874
rect 12544 12850 12572 14486
rect 12728 14482 12756 15438
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13832 15162 13860 15370
rect 13924 15366 13952 16050
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12728 13530 12756 14418
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12912 12986 12940 13738
rect 13004 13326 13032 14758
rect 14292 14414 14320 16050
rect 14752 15910 14780 17614
rect 15304 17202 15332 17614
rect 15396 17270 15424 17614
rect 15856 17338 15884 17614
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 17236 17202 17264 17614
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 17224 17196 17276 17202
rect 17328 17184 17356 17682
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17972 17338 18000 17614
rect 18064 17338 18092 18090
rect 18340 17678 18368 18906
rect 20272 18834 20300 19314
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20364 18970 20392 19246
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 18616 18290 18644 18702
rect 20180 18290 20208 18702
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18248 17270 18276 17546
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 17408 17196 17460 17202
rect 17328 17156 17408 17184
rect 17224 17138 17276 17144
rect 17408 17138 17460 17144
rect 15304 16182 15332 17138
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14476 14958 14504 15846
rect 14752 15570 14780 15846
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14844 15026 14872 15642
rect 15304 15162 15332 16118
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15764 15502 15792 15914
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14384 14618 14412 14894
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 13530 13584 13874
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12636 12442 12664 12718
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 12452 11218 12480 12174
rect 14292 11694 14320 14350
rect 14384 14074 14412 14350
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14476 12442 14504 14894
rect 14936 14618 14964 14894
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14936 13938 14964 14554
rect 15304 14074 15332 15098
rect 15396 14414 15424 15438
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14414 15608 14758
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 15672 13462 15700 15370
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 15660 13456 15712 13462
rect 15660 13398 15712 13404
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14476 11762 14504 12378
rect 15212 11762 15240 13126
rect 15672 12850 15700 13398
rect 16592 13394 16620 14962
rect 17236 13394 17264 17138
rect 18248 15722 18276 17206
rect 18340 17134 18368 17614
rect 20180 17134 20208 18226
rect 20732 17882 20760 18566
rect 20824 18426 20852 18634
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20916 17814 20944 19450
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21008 18290 21036 19110
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21100 18222 21128 19994
rect 21192 19854 21220 20198
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21088 18216 21140 18222
rect 21088 18158 21140 18164
rect 20904 17808 20956 17814
rect 20904 17750 20956 17756
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20352 17604 20404 17610
rect 20352 17546 20404 17552
rect 20364 17338 20392 17546
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20548 17338 20576 17478
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 20640 17202 20668 17682
rect 20916 17202 20944 17750
rect 21088 17672 21140 17678
rect 21192 17660 21220 19790
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21376 18290 21404 19654
rect 21468 19378 21496 20198
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21560 19446 21588 19926
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21548 19440 21600 19446
rect 21548 19382 21600 19388
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21140 17632 21220 17660
rect 21456 17672 21508 17678
rect 21088 17614 21140 17620
rect 21560 17660 21588 19382
rect 21744 18970 21772 19790
rect 21836 19514 21864 20470
rect 23400 20466 23428 21966
rect 22928 20460 22980 20466
rect 22928 20402 22980 20408
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 22008 20324 22060 20330
rect 22008 20266 22060 20272
rect 22020 20058 22048 20266
rect 22560 20256 22612 20262
rect 22560 20198 22612 20204
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 21824 19508 21876 19514
rect 21824 19450 21876 19456
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21744 17678 21772 18906
rect 21836 18290 21864 19450
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 21928 18630 21956 18906
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21928 17678 21956 18566
rect 22020 18290 22048 19314
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22388 18426 22416 19246
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22572 18290 22600 20198
rect 22940 19922 22968 20402
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 22928 19916 22980 19922
rect 22928 19858 22980 19864
rect 22940 19378 22968 19858
rect 23676 19854 23704 19994
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23124 18766 23152 19110
rect 23676 18766 23704 19790
rect 23112 18760 23164 18766
rect 23112 18702 23164 18708
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22664 17746 22692 18022
rect 23676 17746 23704 18702
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 21508 17632 21588 17660
rect 21732 17672 21784 17678
rect 21456 17614 21508 17620
rect 21732 17614 21784 17620
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 21836 17338 21864 17614
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 18156 15694 18276 15722
rect 17408 13796 17460 13802
rect 17408 13738 17460 13744
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 16316 12782 16344 13126
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13464 10810 13492 11018
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 14108 10674 14136 11494
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14384 10538 14412 11698
rect 14476 10674 14504 11698
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14936 11354 14964 11630
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14936 10810 14964 11290
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 15212 10742 15240 11698
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 11082 15884 11494
rect 16040 11354 16068 12038
rect 16316 11762 16344 12038
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16592 11694 16620 13330
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16684 12442 16712 12650
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16776 12306 16804 12582
rect 16868 12442 16896 13262
rect 17132 12844 17184 12850
rect 17236 12832 17264 13330
rect 17184 12804 17264 12832
rect 17132 12786 17184 12792
rect 17236 12714 17264 12804
rect 17420 12782 17448 13738
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17224 12708 17276 12714
rect 17224 12650 17276 12656
rect 17420 12646 17448 12718
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16868 11898 16896 12378
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 17420 11286 17448 12582
rect 17604 11898 17632 13262
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18064 12374 18092 12786
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17880 11762 17908 12106
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17972 11558 18000 12174
rect 18156 11830 18184 15694
rect 20180 14414 20208 17070
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18248 12306 18276 12582
rect 18524 12442 18552 12786
rect 19352 12782 19380 13126
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19444 12714 19472 13262
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 19444 12238 19472 12650
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17972 11354 18000 11494
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 15212 10062 15240 10678
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15948 10062 15976 10406
rect 16224 10130 16252 11086
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17052 10674 17080 10950
rect 18064 10674 18092 11630
rect 18156 11354 18184 11766
rect 19628 11694 19656 14350
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20272 14074 20300 14282
rect 20640 14278 20668 17138
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19996 13258 20024 13738
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19720 12306 19748 13126
rect 19996 12918 20024 13194
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 20088 12782 20116 13262
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 20456 12306 20484 13942
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20548 12986 20576 13874
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20640 12986 20668 13262
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18156 11082 18184 11290
rect 19536 11150 19564 11562
rect 19628 11218 19656 11630
rect 19904 11354 19932 11698
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 20272 11218 20300 12038
rect 20824 11558 20852 13874
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20916 12714 20944 13262
rect 21284 12850 21312 17274
rect 21928 17202 21956 17614
rect 21916 17196 21968 17202
rect 21916 17138 21968 17144
rect 22204 17134 22232 17614
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23124 17202 23152 17478
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22204 16574 22232 17070
rect 23492 16998 23520 17478
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 22848 16658 22876 16934
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 23492 16590 23520 16934
rect 23480 16584 23532 16590
rect 22204 16546 22324 16574
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21652 12850 21680 14214
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20916 12238 20944 12650
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 21180 12096 21232 12102
rect 21284 12084 21312 12786
rect 21744 12782 21772 13330
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21232 12056 21312 12084
rect 21180 12038 21232 12044
rect 21284 11830 21312 12056
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21468 11762 21496 12038
rect 21744 11762 21772 12718
rect 21836 12238 21864 12718
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21836 11898 21864 12174
rect 22296 12170 22324 16546
rect 23480 16526 23532 16532
rect 23676 16454 23704 17138
rect 23768 16574 23796 22066
rect 24320 20058 24348 24074
rect 24504 23882 24532 24142
rect 24504 23854 24624 23882
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24504 23322 24532 23666
rect 24596 23322 24624 23854
rect 24492 23316 24544 23322
rect 24492 23258 24544 23264
rect 24584 23316 24636 23322
rect 24584 23258 24636 23264
rect 24596 22710 24624 23258
rect 24688 23118 24716 24278
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24584 22704 24636 22710
rect 24584 22646 24636 22652
rect 24872 22642 24900 25758
rect 25240 25702 25268 26794
rect 25780 25832 25832 25838
rect 25780 25774 25832 25780
rect 24952 25696 25004 25702
rect 24952 25638 25004 25644
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 24964 24070 24992 25638
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24964 23186 24992 24006
rect 25792 23866 25820 25774
rect 25780 23860 25832 23866
rect 25780 23802 25832 23808
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24492 20392 24544 20398
rect 24492 20334 24544 20340
rect 24308 20052 24360 20058
rect 24308 19994 24360 20000
rect 24320 19514 24348 19994
rect 24308 19508 24360 19514
rect 24308 19450 24360 19456
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23860 18970 23888 19246
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 24504 18834 24532 20334
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 24492 18828 24544 18834
rect 24492 18770 24544 18776
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23860 17542 23888 18566
rect 24044 18290 24072 18770
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 23952 17882 23980 18226
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23952 16590 23980 17682
rect 24044 16658 24072 18226
rect 24688 17678 24716 18838
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24872 17882 24900 18634
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24320 16794 24348 17070
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 23940 16584 23992 16590
rect 23768 16546 23888 16574
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23676 14822 23704 16390
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23216 14074 23244 14282
rect 23204 14068 23256 14074
rect 23204 14010 23256 14016
rect 23676 13326 23704 14758
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22284 12164 22336 12170
rect 22284 12106 22336 12112
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20824 11286 20852 11494
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 21744 11150 21772 11698
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22112 11354 22140 11494
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22204 11150 22232 12038
rect 22296 11354 22324 12106
rect 22480 11898 22508 12786
rect 23032 12782 23060 13126
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23492 12306 23520 12650
rect 23584 12374 23612 12922
rect 23676 12850 23704 13126
rect 23768 12918 23796 13806
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23572 12368 23624 12374
rect 23572 12310 23624 12316
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22756 11898 22784 12174
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 23676 11286 23704 12786
rect 23860 11354 23888 16546
rect 23940 16526 23992 16532
rect 23952 15910 23980 16526
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 23952 13190 23980 15846
rect 24044 14906 24072 16594
rect 24964 16590 24992 16934
rect 27540 16794 27568 17138
rect 28264 17128 28316 17134
rect 28262 17096 28264 17105
rect 28316 17096 28318 17105
rect 28262 17031 28318 17040
rect 27528 16788 27580 16794
rect 27528 16730 27580 16736
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 27080 16114 27108 16390
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 28264 16040 28316 16046
rect 28264 15982 28316 15988
rect 28276 15745 28304 15982
rect 28262 15736 28318 15745
rect 28262 15671 28318 15680
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 24044 14878 24164 14906
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 23940 13184 23992 13190
rect 23940 13126 23992 13132
rect 24044 12850 24072 14758
rect 24136 14414 24164 14878
rect 25148 14618 25176 14962
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 25424 14618 25452 14894
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 24860 14408 24912 14414
rect 28448 14408 28500 14414
rect 24860 14350 24912 14356
rect 28446 14376 28448 14385
rect 28500 14376 28502 14385
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24136 11762 24164 14350
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24228 12918 24256 13670
rect 24412 13462 24440 13806
rect 24400 13456 24452 13462
rect 24400 13398 24452 13404
rect 24872 12986 24900 14350
rect 28446 14311 28502 14320
rect 24952 13932 25004 13938
rect 24952 13874 25004 13880
rect 24964 12986 24992 13874
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 24492 11688 24544 11694
rect 24492 11630 24544 11636
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23664 11280 23716 11286
rect 23664 11222 23716 11228
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18248 10810 18276 11086
rect 19536 10810 19564 11086
rect 23860 11082 23888 11290
rect 24504 11150 24532 11630
rect 24596 11558 24624 12786
rect 24780 11898 24808 12786
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 25148 11762 25176 12038
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24780 11286 24808 11630
rect 24768 11280 24820 11286
rect 24768 11222 24820 11228
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 28264 11076 28316 11082
rect 28264 11018 28316 11024
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18064 10266 18092 10610
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15764 9722 15792 9998
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 28276 8634 28304 11018
rect 28264 8628 28316 8634
rect 28264 8570 28316 8576
rect 28276 8090 28304 8570
rect 28448 8492 28500 8498
rect 28448 8434 28500 8440
rect 28460 8265 28488 8434
rect 28446 8256 28502 8265
rect 28446 8191 28502 8200
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5828 800 5856 2382
rect 21928 800 21956 2382
rect 5814 0 5870 800
rect 21914 0 21970 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 110 44512 166 44568
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 1214 38120 1270 38176
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 846 32172 848 32192
rect 848 32172 900 32192
rect 900 32172 902 32192
rect 846 32136 902 32172
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 1306 29960 1362 30016
rect 846 29416 902 29472
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 846 23976 902 24032
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 846 23296 902 23352
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 1214 21800 1270 21856
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 846 17856 902 17912
rect 1306 17040 1362 17096
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 28262 32000 28318 32056
rect 28446 31320 28502 31376
rect 28446 27240 28502 27296
rect 28262 17076 28264 17096
rect 28264 17076 28316 17096
rect 28316 17076 28318 17096
rect 28262 17040 28318 17076
rect 28262 15680 28318 15736
rect 28446 14356 28448 14376
rect 28448 14356 28500 14376
rect 28500 14356 28502 14376
rect 28446 14320 28502 14356
rect 28446 8200 28502 8256
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 105 44570 171 44573
rect 105 44568 1042 44570
rect 105 44512 110 44568
rect 166 44512 1042 44568
rect 105 44510 1042 44512
rect 105 44507 171 44510
rect 0 44298 800 44328
rect 982 44298 1042 44510
rect 0 44238 1042 44298
rect 0 44208 800 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 0 38178 800 38208
rect 1209 38178 1275 38181
rect 0 38176 1275 38178
rect 0 38120 1214 38176
rect 1270 38120 1275 38176
rect 0 38118 1275 38120
rect 0 38088 800 38118
rect 1209 38115 1275 38118
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 841 32194 907 32197
rect 798 32192 907 32194
rect 798 32136 846 32192
rect 902 32136 907 32192
rect 798 32131 907 32136
rect 798 32088 858 32131
rect 0 31998 858 32088
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 28257 32058 28323 32061
rect 29200 32058 30000 32088
rect 28257 32056 30000 32058
rect 28257 32000 28262 32056
rect 28318 32000 30000 32056
rect 28257 31998 30000 32000
rect 0 31968 800 31998
rect 28257 31995 28323 31998
rect 29200 31968 30000 31998
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 28441 31378 28507 31381
rect 29200 31378 30000 31408
rect 28441 31376 30000 31378
rect 28441 31320 28446 31376
rect 28502 31320 30000 31376
rect 28441 31318 30000 31320
rect 28441 31315 28507 31318
rect 29200 31288 30000 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 0 30018 800 30048
rect 1301 30018 1367 30021
rect 0 30016 1367 30018
rect 0 29960 1306 30016
rect 1362 29960 1367 30016
rect 0 29958 1367 29960
rect 0 29928 800 29958
rect 1301 29955 1367 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 841 29474 907 29477
rect 798 29472 907 29474
rect 798 29416 846 29472
rect 902 29416 907 29472
rect 798 29411 907 29416
rect 798 29368 858 29411
rect 0 29278 858 29368
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 0 29248 800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 28441 27298 28507 27301
rect 29200 27298 30000 27328
rect 28441 27296 30000 27298
rect 28441 27240 28446 27296
rect 28502 27240 30000 27296
rect 28441 27238 30000 27240
rect 28441 27235 28507 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 29200 27208 30000 27238
rect 4870 27167 5186 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 841 24034 907 24037
rect 798 24032 907 24034
rect 798 23976 846 24032
rect 902 23976 907 24032
rect 798 23971 907 23976
rect 798 23928 858 23971
rect 0 23838 858 23928
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 0 23808 800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 841 23354 907 23357
rect 798 23352 907 23354
rect 798 23296 846 23352
rect 902 23296 907 23352
rect 798 23291 907 23296
rect 798 23248 858 23291
rect 0 23158 858 23248
rect 0 23128 800 23158
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 0 21858 800 21888
rect 1209 21858 1275 21861
rect 0 21856 1275 21858
rect 0 21800 1214 21856
rect 1270 21800 1275 21856
rect 0 21798 1275 21800
rect 0 21768 800 21798
rect 1209 21795 1275 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 841 17914 907 17917
rect 798 17912 907 17914
rect 798 17856 846 17912
rect 902 17856 907 17912
rect 798 17851 907 17856
rect 798 17808 858 17851
rect 0 17718 858 17808
rect 0 17688 800 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 0 17098 800 17128
rect 1301 17098 1367 17101
rect 0 17096 1367 17098
rect 0 17040 1306 17096
rect 1362 17040 1367 17096
rect 0 17038 1367 17040
rect 0 17008 800 17038
rect 1301 17035 1367 17038
rect 28257 17098 28323 17101
rect 29200 17098 30000 17128
rect 28257 17096 30000 17098
rect 28257 17040 28262 17096
rect 28318 17040 30000 17096
rect 28257 17038 30000 17040
rect 28257 17035 28323 17038
rect 29200 17008 30000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 28257 15738 28323 15741
rect 29200 15738 30000 15768
rect 28257 15736 30000 15738
rect 28257 15680 28262 15736
rect 28318 15680 30000 15736
rect 28257 15678 30000 15680
rect 28257 15675 28323 15678
rect 29200 15648 30000 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 28441 14378 28507 14381
rect 29200 14378 30000 14408
rect 28441 14376 30000 14378
rect 28441 14320 28446 14376
rect 28502 14320 30000 14376
rect 28441 14318 30000 14320
rect 28441 14315 28507 14318
rect 29200 14288 30000 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 28441 8258 28507 8261
rect 29200 8258 30000 8288
rect 28441 8256 30000 8258
rect 28441 8200 28446 8256
rect 28502 8200 30000 8256
rect 28441 8198 30000 8200
rect 28441 8195 28507 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 29200 8168 30000 8198
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 46816 5188 47376
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1
transform -1 0 23828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1
transform -1 0 22632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1
transform -1 0 21528 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1
transform -1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1
transform 1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1
transform -1 0 14904 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1
transform 1 0 14628 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1
transform -1 0 25760 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1
transform -1 0 25024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1
transform -1 0 23828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1
transform 1 0 21344 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1
transform -1 0 20056 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1
transform -1 0 19596 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1
transform -1 0 16468 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1
transform 1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1
transform -1 0 16100 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1
transform 1 0 12512 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1
transform 1 0 13524 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1
transform -1 0 13064 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1
transform 1 0 14168 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1
transform -1 0 13616 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _382_
timestamp 1
transform -1 0 9476 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _383_
timestamp 1
transform 1 0 6624 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _384_
timestamp 1
transform -1 0 8280 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _385_
timestamp 1
transform 1 0 7268 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _386_
timestamp 1
transform 1 0 7360 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _387_
timestamp 1
transform -1 0 6072 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _388_
timestamp 1
transform -1 0 8188 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _389_
timestamp 1
transform 1 0 7820 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _390_
timestamp 1
transform -1 0 11224 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _391_
timestamp 1
transform -1 0 4968 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _392_
timestamp 1
transform -1 0 5888 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _393_
timestamp 1
transform -1 0 6348 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _394_
timestamp 1
transform 1 0 9016 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _395_
timestamp 1
transform 1 0 6532 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _396_
timestamp 1
transform -1 0 9476 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _397_
timestamp 1
transform -1 0 5428 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _398_
timestamp 1
transform 1 0 6440 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _399_
timestamp 1
transform -1 0 5336 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _400_
timestamp 1
transform 1 0 4784 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _401_
timestamp 1
transform 1 0 6440 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _402_
timestamp 1
transform 1 0 6440 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _403_
timestamp 1
transform 1 0 5428 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _404_
timestamp 1
transform 1 0 5612 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _405_
timestamp 1
transform 1 0 2484 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _406_
timestamp 1
transform -1 0 5520 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _407_
timestamp 1
transform 1 0 4140 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _408_
timestamp 1
transform 1 0 5520 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _409_
timestamp 1
transform -1 0 8372 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _410_
timestamp 1
transform -1 0 13156 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _411_
timestamp 1
transform 1 0 11592 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _412_
timestamp 1
transform -1 0 13064 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _413_
timestamp 1
transform 1 0 11408 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _414_
timestamp 1
transform -1 0 14720 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _415_
timestamp 1
transform -1 0 12788 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _416_
timestamp 1
transform -1 0 11132 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _417_
timestamp 1
transform -1 0 10764 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _418_
timestamp 1
transform -1 0 13800 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _419_
timestamp 1
transform 1 0 4232 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _420_
timestamp 1
transform 1 0 8280 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _421_
timestamp 1
transform -1 0 11132 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _422_
timestamp 1
transform 1 0 12052 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _423_
timestamp 1
transform 1 0 13248 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _424_
timestamp 1
transform -1 0 12512 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _425_
timestamp 1
transform -1 0 8556 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _426_
timestamp 1
transform 1 0 8280 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _427_
timestamp 1
transform 1 0 7912 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _428_
timestamp 1
transform 1 0 9016 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _429_
timestamp 1
transform -1 0 10672 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _430_
timestamp 1
transform -1 0 8740 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _431_
timestamp 1
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _432_
timestamp 1
transform 1 0 10488 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _433_
timestamp 1
transform 1 0 3588 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _434_
timestamp 1
transform -1 0 6900 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _435_
timestamp 1
transform -1 0 11316 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _436_
timestamp 1
transform -1 0 8004 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _437_
timestamp 1
transform -1 0 9476 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _438_
timestamp 1
transform -1 0 12052 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _439_
timestamp 1
transform -1 0 8372 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _440_
timestamp 1
transform 1 0 9016 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _441_
timestamp 1
transform 1 0 9016 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _442_
timestamp 1
transform 1 0 6624 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _443_
timestamp 1
transform -1 0 10396 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _444_
timestamp 1
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _445_
timestamp 1
transform 1 0 12512 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _446_
timestamp 1
transform -1 0 10212 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _447_
timestamp 1
transform 1 0 5428 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _448_
timestamp 1
transform -1 0 6164 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _449_
timestamp 1
transform -1 0 8004 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _450_
timestamp 1
transform -1 0 9936 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _451_
timestamp 1
transform 1 0 10212 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _452_
timestamp 1
transform -1 0 9752 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _453_
timestamp 1
transform -1 0 7544 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _454_
timestamp 1
transform 1 0 7728 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _455_
timestamp 1
transform -1 0 5888 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _456_
timestamp 1
transform 1 0 10396 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _457_
timestamp 1
transform 1 0 6900 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _458_
timestamp 1
transform -1 0 11500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _459_
timestamp 1
transform -1 0 6992 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _460_
timestamp 1
transform 1 0 9016 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _461_
timestamp 1
transform 1 0 14904 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _462_
timestamp 1
transform 1 0 16192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _463_
timestamp 1
transform 1 0 14996 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _464_
timestamp 1
transform -1 0 15824 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _465_
timestamp 1
transform -1 0 16468 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _466_
timestamp 1
transform -1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _467_
timestamp 1
transform -1 0 19044 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _468_
timestamp 1
transform -1 0 18400 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _469_
timestamp 1
transform 1 0 17388 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _470_
timestamp 1
transform 1 0 19780 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _471_
timestamp 1
transform 1 0 20976 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _472_
timestamp 1
transform -1 0 19872 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _473_
timestamp 1
transform 1 0 21068 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _474_
timestamp 1
transform 1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _475_
timestamp 1
transform 1 0 20792 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _476_
timestamp 1
transform 1 0 21896 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _477_
timestamp 1
transform 1 0 22540 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _478_
timestamp 1
transform -1 0 22448 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _479_
timestamp 1
transform 1 0 23644 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _480_
timestamp 1
transform 1 0 24472 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _481_
timestamp 1
transform 1 0 2944 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _482_
timestamp 1
transform 1 0 4048 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _483_
timestamp 1
transform 1 0 5060 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _484_
timestamp 1
transform 1 0 5704 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _485_
timestamp 1
transform 1 0 5980 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _486_
timestamp 1
transform 1 0 9016 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _487_
timestamp 1
transform 1 0 10488 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _488_
timestamp 1
transform 1 0 9844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _489_
timestamp 1
transform 1 0 10672 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _490_
timestamp 1
transform -1 0 14536 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _491_
timestamp 1
transform 1 0 14260 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _492_
timestamp 1
transform 1 0 9660 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _493_
timestamp 1
transform -1 0 10304 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _494_
timestamp 1
transform 1 0 12052 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _495_
timestamp 1
transform -1 0 11316 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _496_
timestamp 1
transform 1 0 11592 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _497_
timestamp 1
transform 1 0 11684 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _498_
timestamp 1
transform 1 0 11592 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _499_
timestamp 1
transform 1 0 12604 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _500_
timestamp 1
transform 1 0 12236 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _501_
timestamp 1
transform 1 0 11684 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _502_
timestamp 1
transform -1 0 13156 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _503_
timestamp 1
transform -1 0 11316 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _504_
timestamp 1
transform -1 0 12512 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _505_
timestamp 1
transform 1 0 10948 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _506_
timestamp 1
transform -1 0 12328 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _507_
timestamp 1
transform 1 0 10304 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _508_
timestamp 1
transform -1 0 12236 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _509_
timestamp 1
transform 1 0 10764 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _510_
timestamp 1
transform 1 0 13892 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _511_
timestamp 1
transform -1 0 13524 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _512_
timestamp 1
transform -1 0 12696 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _513_
timestamp 1
transform -1 0 11408 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _514_
timestamp 1
transform 1 0 9200 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _515_
timestamp 1
transform 1 0 13156 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _516_
timestamp 1
transform 1 0 11592 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _517_
timestamp 1
transform -1 0 14352 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _518_
timestamp 1
transform -1 0 12052 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _519_
timestamp 1
transform 1 0 10396 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _520_
timestamp 1
transform 1 0 11500 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _521_
timestamp 1
transform -1 0 12236 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _522_
timestamp 1
transform 1 0 9844 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _523_
timestamp 1
transform 1 0 10488 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _524_
timestamp 1
transform 1 0 9384 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _525_
timestamp 1
transform 1 0 10488 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _526_
timestamp 1
transform -1 0 14076 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _527_
timestamp 1
transform -1 0 13616 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _528_
timestamp 1
transform -1 0 13892 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _529_
timestamp 1
transform -1 0 12972 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _530_
timestamp 1
transform 1 0 11592 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _531_
timestamp 1
transform 1 0 13248 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _532_
timestamp 1
transform 1 0 14628 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _533_
timestamp 1
transform -1 0 14720 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _534_
timestamp 1
transform -1 0 13064 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _535_
timestamp 1
transform -1 0 14812 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _536_
timestamp 1
transform 1 0 13800 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _537_
timestamp 1
transform 1 0 14168 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _538_
timestamp 1
transform 1 0 14628 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _539_
timestamp 1
transform 1 0 13248 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _540_
timestamp 1
transform 1 0 14168 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _541_
timestamp 1
transform -1 0 13984 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _542_
timestamp 1
transform 1 0 14168 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _543_
timestamp 1
transform -1 0 16008 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _544_
timestamp 1
transform 1 0 16284 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_2  _545_
timestamp 1
transform -1 0 15272 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_2  _546_
timestamp 1
transform 1 0 13248 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _547_
timestamp 1
transform 1 0 16744 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _548_
timestamp 1
transform -1 0 18216 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _549_
timestamp 1
transform -1 0 17388 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _550_
timestamp 1
transform -1 0 17940 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _551_
timestamp 1
transform 1 0 16744 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _552_
timestamp 1
transform 1 0 15640 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _553_
timestamp 1
transform 1 0 16468 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _554_
timestamp 1
transform -1 0 15364 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _555_
timestamp 1
transform -1 0 17940 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _556_
timestamp 1
transform -1 0 18952 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _557_
timestamp 1
transform -1 0 19044 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _558_
timestamp 1
transform -1 0 18032 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _559_
timestamp 1
transform 1 0 18216 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _560_
timestamp 1
transform 1 0 19320 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _561_
timestamp 1
transform -1 0 17572 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _562_
timestamp 1
transform 1 0 18584 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _563_
timestamp 1
transform -1 0 18860 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _564_
timestamp 1
transform -1 0 19596 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _565_
timestamp 1
transform 1 0 17480 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _566_
timestamp 1
transform 1 0 19412 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _567_
timestamp 1
transform 1 0 17480 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _568_
timestamp 1
transform 1 0 20516 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _569_
timestamp 1
transform 1 0 21896 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _570_
timestamp 1
transform -1 0 23000 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _571_
timestamp 1
transform 1 0 18676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _572_
timestamp 1
transform -1 0 19964 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _573_
timestamp 1
transform 1 0 20976 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _574_
timestamp 1
transform 1 0 21160 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _575_
timestamp 1
transform 1 0 20884 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _576_
timestamp 1
transform -1 0 22540 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _577_
timestamp 1
transform 1 0 20976 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _578_
timestamp 1
transform 1 0 20884 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _579_
timestamp 1
transform 1 0 21712 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _580_
timestamp 1
transform -1 0 21620 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _581_
timestamp 1
transform 1 0 23736 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _582_
timestamp 1
transform 1 0 22908 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _583_
timestamp 1
transform -1 0 24932 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _584_
timestamp 1
transform 1 0 22724 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _585_
timestamp 1
transform -1 0 22356 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _586_
timestamp 1
transform 1 0 23552 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _587_
timestamp 1
transform -1 0 24564 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _588_
timestamp 1
transform -1 0 23552 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _589_
timestamp 1
transform -1 0 24288 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _590_
timestamp 1
transform -1 0 26036 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _591_
timestamp 1
transform -1 0 24840 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _592_
timestamp 1
transform 1 0 25024 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _593_
timestamp 1
transform -1 0 24012 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _594_
timestamp 1
transform 1 0 11592 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _595_
timestamp 1
transform 1 0 13064 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _596_
timestamp 1
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _597_
timestamp 1
transform 1 0 12420 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _598_
timestamp 1
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _599_
timestamp 1
transform 1 0 14168 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_2  _600_
timestamp 1
transform 1 0 11776 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_2  _601_
timestamp 1
transform 1 0 12328 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _602_
timestamp 1
transform -1 0 14996 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _603_
timestamp 1
transform 1 0 14904 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _604_
timestamp 1
transform -1 0 14444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _605_
timestamp 1
transform 1 0 13432 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _606_
timestamp 1
transform 1 0 15364 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _607_
timestamp 1
transform 1 0 13064 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _608_
timestamp 1
transform 1 0 13892 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _609_
timestamp 1
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _610_
timestamp 1
transform 1 0 15180 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _611_
timestamp 1
transform -1 0 19044 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _612_
timestamp 1
transform -1 0 16928 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _613_
timestamp 1
transform 1 0 15824 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _614_
timestamp 1
transform 1 0 16744 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _615_
timestamp 1
transform -1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _616_
timestamp 1
transform -1 0 18308 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _617_
timestamp 1
transform -1 0 17388 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _618_
timestamp 1
transform 1 0 15456 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _619_
timestamp 1
transform 1 0 17020 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _620_
timestamp 1
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _621_
timestamp 1
transform -1 0 20700 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _622_
timestamp 1
transform 1 0 17572 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _623_
timestamp 1
transform 1 0 17112 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _624_
timestamp 1
transform 1 0 19228 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _625_
timestamp 1
transform -1 0 20884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _626_
timestamp 1
transform -1 0 19412 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _627_
timestamp 1
transform -1 0 21528 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _628_
timestamp 1
transform -1 0 20332 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _629_
timestamp 1
transform 1 0 19412 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _630_
timestamp 1
transform 1 0 20240 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _631_
timestamp 1
transform -1 0 19964 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _632_
timestamp 1
transform 1 0 24472 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _633_
timestamp 1
transform 1 0 21712 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _634_
timestamp 1
transform 1 0 21988 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _635_
timestamp 1
transform -1 0 22448 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _636_
timestamp 1
transform -1 0 21160 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _637_
timestamp 1
transform 1 0 22908 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _638_
timestamp 1
transform -1 0 23920 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _639_
timestamp 1
transform 1 0 25116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _640_
timestamp 1
transform -1 0 25024 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _641_
timestamp 1
transform 1 0 23000 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _642_
timestamp 1
transform -1 0 24748 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _643_
timestamp 1
transform 1 0 25392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _644_
timestamp 1
transform -1 0 24288 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _645_
timestamp 1
transform 1 0 16008 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _646_
timestamp 1
transform 1 0 15824 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _647_
timestamp 1
transform -1 0 14720 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _648_
timestamp 1
transform 1 0 15548 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _649_
timestamp 1
transform -1 0 16192 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _650_
timestamp 1
transform -1 0 16100 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _651_
timestamp 1
transform -1 0 15732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _652_
timestamp 1
transform 1 0 14444 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _653_
timestamp 1
transform 1 0 14168 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _654_
timestamp 1
transform 1 0 14628 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _655_
timestamp 1
transform 1 0 15364 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _656_
timestamp 1
transform 1 0 16100 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _657_
timestamp 1
transform 1 0 16744 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _658_
timestamp 1
transform 1 0 16652 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _659_
timestamp 1
transform -1 0 17940 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _660_
timestamp 1
transform 1 0 22264 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _661_
timestamp 1
transform -1 0 17756 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _662_
timestamp 1
transform 1 0 17940 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _663_
timestamp 1
transform -1 0 19412 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _664_
timestamp 1
transform -1 0 18860 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _665_
timestamp 1
transform 1 0 19872 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _666_
timestamp 1
transform 1 0 21896 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _667_
timestamp 1
transform 1 0 22816 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _668_
timestamp 1
transform 1 0 23736 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_1  _669_
timestamp 1
transform -1 0 25300 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _670_
timestamp 1
transform 1 0 14444 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _671_
timestamp 1
transform 1 0 16008 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _672_
timestamp 1
transform -1 0 15364 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _673_
timestamp 1
transform -1 0 16008 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _674_
timestamp 1
transform 1 0 16744 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _675_
timestamp 1
transform -1 0 16468 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _676_
timestamp 1
transform -1 0 19964 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _677_
timestamp 1
transform 1 0 19504 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _678_
timestamp 1
transform -1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _679_
timestamp 1
transform 1 0 16928 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _680_
timestamp 1
transform 1 0 19964 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _681_
timestamp 1
transform -1 0 18952 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _682_
timestamp 1
transform 1 0 17572 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _683_
timestamp 1
transform 1 0 19320 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _684_
timestamp 1
transform -1 0 18952 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _685_
timestamp 1
transform 1 0 20056 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _686_
timestamp 1
transform 1 0 20700 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _687_
timestamp 1
transform 1 0 19320 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _688_
timestamp 1
transform 1 0 20332 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _689_
timestamp 1
transform -1 0 17572 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _690_
timestamp 1
transform 1 0 22172 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _691_
timestamp 1
transform -1 0 20884 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _692_
timestamp 1
transform -1 0 15640 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _693_
timestamp 1
transform 1 0 15456 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _694_
timestamp 1
transform 1 0 15916 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _695_
timestamp 1
transform -1 0 17664 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _696_
timestamp 1
transform -1 0 19872 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _697_
timestamp 1
transform 1 0 17848 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _698_
timestamp 1
transform 1 0 20148 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _699_
timestamp 1
transform 1 0 21528 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _700_
timestamp 1
transform 1 0 22816 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _701_
timestamp 1
transform 1 0 23460 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _702_
timestamp 1
transform 1 0 15640 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _703_
timestamp 1
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _704_
timestamp 1
transform 1 0 17296 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _705_
timestamp 1
transform -1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _706_
timestamp 1
transform 1 0 18032 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _707_
timestamp 1
transform -1 0 18584 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _708_
timestamp 1
transform -1 0 20240 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _709_
timestamp 1
transform 1 0 19780 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _710_
timestamp 1
transform 1 0 19320 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _711_
timestamp 1
transform 1 0 20884 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _712_
timestamp 1
transform -1 0 21252 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _713_
timestamp 1
transform -1 0 20700 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _714_
timestamp 1
transform -1 0 24012 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _715_
timestamp 1
transform 1 0 23092 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _716_
timestamp 1
transform 1 0 21896 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _717_
timestamp 1
transform 1 0 23368 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _718_
timestamp 1
transform 1 0 24012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _719_
timestamp 1
transform 1 0 22632 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _720_
timestamp 1
transform -1 0 24840 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _721_
timestamp 1
transform 1 0 24472 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _722_
timestamp 1
transform 1 0 8372 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _723_
timestamp 1
transform 1 0 4416 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _724_
timestamp 1
transform 1 0 5060 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _725_
timestamp 1
transform 1 0 4692 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _726_
timestamp 1
transform 1 0 5612 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _727_
timestamp 1
transform 1 0 7912 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _728_
timestamp 1
transform 1 0 9568 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _729_
timestamp 1
transform -1 0 8556 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _730_
timestamp 1
transform 1 0 7176 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _731_
timestamp 1
transform 1 0 7268 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _732_
timestamp 1
transform 1 0 3128 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _733_
timestamp 1
transform 1 0 4968 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _734_
timestamp 1
transform -1 0 7912 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _735_
timestamp 1
transform 1 0 5244 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _736_
timestamp 1
transform 1 0 4232 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _737_
timestamp 1
transform 1 0 5336 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _738_
timestamp 1
transform -1 0 6992 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _739_
timestamp 1
transform -1 0 7912 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _740_
timestamp 1
transform 1 0 12144 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _741_
timestamp 1
transform 1 0 5612 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _742_
timestamp 1
transform 1 0 8648 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _743_
timestamp 1
transform -1 0 10672 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _744_
timestamp 1
transform 1 0 9384 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _745_
timestamp 1
transform 1 0 10488 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _746_
timestamp 1
transform 1 0 12144 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _747_
timestamp 1
transform -1 0 13892 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _748_
timestamp 1
transform -1 0 14076 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _749_
timestamp 1
transform 1 0 11592 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _750_
timestamp 1
transform 1 0 4508 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _751_
timestamp 1
transform 1 0 6440 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _752_
timestamp 1
transform 1 0 9844 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _753_
timestamp 1
transform -1 0 11316 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _754_
timestamp 1
transform -1 0 10488 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _755_
timestamp 1
transform 1 0 7176 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _756_
timestamp 1
transform 1 0 6992 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _757_
timestamp 1
transform 1 0 8648 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _758_
timestamp 1
transform 1 0 10580 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _759_
timestamp 1
transform 1 0 5428 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _760_
timestamp 1
transform 1 0 5612 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _761_
timestamp 1
transform 1 0 6716 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _762_
timestamp 1
transform 1 0 7268 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _763_
timestamp 1
transform 1 0 9936 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _764_
timestamp 1
transform -1 0 10028 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _765_
timestamp 1
transform 1 0 7268 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _766_
timestamp 1
transform -1 0 13064 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _767_
timestamp 1
transform 1 0 9752 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _768_
timestamp 1
transform 1 0 14536 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _769_
timestamp 1
transform 1 0 14536 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _770_
timestamp 1
transform 1 0 15916 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _771_
timestamp 1
transform 1 0 17572 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _772_
timestamp 1
transform 1 0 18124 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _773_
timestamp 1
transform 1 0 20332 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _774_
timestamp 1
transform -1 0 23460 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _775_
timestamp 1
transform -1 0 24104 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _776_
timestamp 1
transform 1 0 8924 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _777_
timestamp 1
transform 1 0 3312 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _778_
timestamp 1
transform 1 0 4600 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _779_
timestamp 1
transform 1 0 4692 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _780_
timestamp 1
transform 1 0 5244 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _781_
timestamp 1
transform 1 0 6808 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _782_
timestamp 1
transform 1 0 8096 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _783_
timestamp 1
transform -1 0 9292 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _784_
timestamp 1
transform 1 0 6440 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _785_
timestamp 1
transform -1 0 13892 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _786_
timestamp 1
transform 1 0 12420 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _787_
timestamp 1
transform -1 0 12512 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _788_
timestamp 1
transform 1 0 14168 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _789_
timestamp 1
transform 1 0 9844 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _790_
timestamp 1
transform 1 0 9844 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _791_
timestamp 1
transform 1 0 14168 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _792_
timestamp 1
transform 1 0 14996 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _793_
timestamp 1
transform 1 0 12420 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _794_
timestamp 1
transform 1 0 9016 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _795_
timestamp 1
transform 1 0 14996 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _796_
timestamp 1
transform 1 0 14812 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _797_
timestamp 1
transform 1 0 17572 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _798_
timestamp 1
transform 1 0 17756 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _799_
timestamp 1
transform 1 0 20792 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _800_
timestamp 1
transform 1 0 21896 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _801_
timestamp 1
transform 1 0 22724 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _802_
timestamp 1
transform 1 0 24104 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _803_
timestamp 1
transform 1 0 10672 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _804_
timestamp 1
transform 1 0 12052 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _805_
timestamp 1
transform 1 0 12420 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _806_
timestamp 1
transform 1 0 12972 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _807_
timestamp 1
transform 1 0 15364 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _808_
timestamp 1
transform 1 0 16192 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _809_
timestamp 1
transform -1 0 20792 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _810_
timestamp 1
transform 1 0 19596 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp 1
transform -1 0 24196 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _812_
timestamp 1
transform 1 0 22724 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp 1
transform 1 0 19412 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _814_
timestamp 1
transform 1 0 9936 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _815_
timestamp 1
transform 1 0 25300 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _816_
timestamp 1
transform 1 0 14996 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _817_
timestamp 1
transform 1 0 14904 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _818_
timestamp 1
transform -1 0 17664 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _819_
timestamp 1
transform 1 0 17572 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _820_
timestamp 1
transform -1 0 19320 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _821_
timestamp 1
transform 1 0 18216 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _822_
timestamp 1
transform 1 0 17756 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _823_
timestamp 1
transform 1 0 17112 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _824_
timestamp 1
transform 1 0 24656 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _825_
timestamp 1
transform 1 0 15548 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _826_
timestamp 1
transform 1 0 16744 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _827_
timestamp 1
transform -1 0 19872 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _828_
timestamp 1
transform 1 0 19320 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _829_
timestamp 1
transform -1 0 21528 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _830_
timestamp 1
transform 1 0 21436 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _831_
timestamp 1
transform 1 0 22356 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _832_
timestamp 1
transform 1 0 23828 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _843_
timestamp 1
transform -1 0 27784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__B
timestamp 1
transform -1 0 8648 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__B
timestamp 1
transform 1 0 9660 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__B
timestamp 1
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__B
timestamp 1
transform 1 0 7176 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__B
timestamp 1
transform 1 0 5520 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__B
timestamp 1
transform 1 0 4876 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__B
timestamp 1
transform 1 0 3772 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__B
timestamp 1
transform 1 0 5152 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__B
timestamp 1
transform 1 0 8556 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__B
timestamp 1
transform 1 0 12328 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__B
timestamp 1
transform -1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__B
timestamp 1
transform 1 0 10304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__B
timestamp 1
transform 1 0 10948 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1
transform 1 0 4876 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__B
timestamp 1
transform 1 0 8924 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__B
timestamp 1
transform 1 0 11132 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__B
timestamp 1
transform 1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__B
timestamp 1
transform 1 0 13892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__B
timestamp 1
transform -1 0 12880 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__B
timestamp 1
transform 1 0 8556 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__B
timestamp 1
transform 1 0 8740 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__B
timestamp 1
transform 1 0 7544 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1
transform 1 0 4232 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__B
timestamp 1
transform 1 0 5980 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__B
timestamp 1
transform 1 0 11500 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__B
timestamp 1
transform -1 0 7360 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__B
timestamp 1
transform 1 0 9660 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__B
timestamp 1
transform 1 0 8372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__B1
timestamp 1
transform 1 0 24196 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__B
timestamp 1
transform 1 0 5612 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__B1
timestamp 1
transform 1 0 14720 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__C1
timestamp 1
transform 1 0 12972 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__C1
timestamp 1
transform -1 0 13892 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__A
timestamp 1
transform 1 0 14904 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__538__C1
timestamp 1
transform 1 0 15364 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__B1
timestamp 1
transform 1 0 16192 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A
timestamp 1
transform 1 0 15364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__A
timestamp 1
transform 1 0 17572 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__C1
timestamp 1
transform 1 0 18032 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__A
timestamp 1
transform -1 0 20700 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__A
timestamp 1
transform 1 0 20976 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__588__A
timestamp 1
transform -1 0 25392 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__593__C1
timestamp 1
transform 1 0 24012 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__598__B1
timestamp 1
transform 1 0 14904 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__A
timestamp 1
transform 1 0 14168 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__615__A
timestamp 1
transform 1 0 16100 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__A
timestamp 1
transform -1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__B1
timestamp 1
transform 1 0 21068 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__A
timestamp 1
transform 1 0 19964 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__A
timestamp 1
transform 1 0 25576 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__C1
timestamp 1
transform 1 0 23828 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__659__B1
timestamp 1
transform 1 0 17940 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__670__B
timestamp 1
transform 1 0 14720 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__671__B1
timestamp 1
transform 1 0 16744 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__A
timestamp 1
transform 1 0 16468 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__677__A
timestamp 1
transform 1 0 20424 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__680__A
timestamp 1
transform 1 0 20792 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__683__A
timestamp 1
transform 1 0 19780 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__686__A
timestamp 1
transform 1 0 21160 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__688__B1
timestamp 1
transform 1 0 20884 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__701__B1
timestamp 1
transform 1 0 24012 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__720__B1
timestamp 1
transform -1 0 25208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__843__A
timestamp 1
transform -1 0 28152 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1
transform -1 0 14352 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 1
transform 1 0 16100 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_clk_A
timestamp 1
transform 1 0 11316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_clk_A
timestamp 1
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_clk_A
timestamp 1
transform 1 0 18032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_clk_A
timestamp 1
transform 1 0 16836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_clk_A
timestamp 1
transform 1 0 9108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_clk_A
timestamp 1
transform 1 0 9016 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_clk_A
timestamp 1
transform 1 0 16928 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_clk_A
timestamp 1
transform -1 0 16468 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout12_A
timestamp 1
transform 1 0 12144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout13_X
timestamp 1
transform 1 0 13064 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout14_X
timestamp 1
transform 1 0 13248 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout16_A
timestamp 1
transform 1 0 23460 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout17_A
timestamp 1
transform 1 0 23828 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout17_X
timestamp 1
transform 1 0 24472 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout18_A
timestamp 1
transform 1 0 23184 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout18_X
timestamp 1
transform 1 0 24472 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1
transform -1 0 5888 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1
transform -1 0 2116 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1
transform -1 0 2116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1
transform -1 0 2116 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1
transform -1 0 6624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1
transform -1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1
transform -1 0 27968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_X
timestamp 1
transform -1 0 28520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform 1 0 14076 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1
transform -1 0 11132 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1
transform 1 0 8096 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1
transform 1 0 18400 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1
transform 1 0 17204 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1
transform 1 0 7084 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1
transform -1 0 8740 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1
transform 1 0 16744 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1
transform 1 0 16376 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinvlp_4  clkload0
timestamp 1
transform 1 0 9292 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload1
timestamp 1
transform 1 0 7728 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_16  clkload2
timestamp 1
transform 1 0 18400 0 -1 18496
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_8  clkload3
timestamp 1
transform 1 0 7084 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  clkload4
timestamp 1
transform 1 0 6900 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload5
timestamp 1
transform 1 0 16744 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  clkload6
timestamp 1
transform 1 0 16744 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  fanout12
timestamp 1
transform -1 0 11960 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1
transform -1 0 12880 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1
transform 1 0 12512 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout15
timestamp 1
transform 1 0 13524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout16
timestamp 1
transform 1 0 22724 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1
transform 1 0 23092 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout18
timestamp 1
transform 1 0 23552 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_3
timestamp 1562078211
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_15
timestamp 1562078211
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_29
timestamp 1562078211
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_0_41
timestamp 1
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51
timestamp 1
transform 1 0 5796 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_60
timestamp 1562078211
transform 1 0 6624 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_72
timestamp 1562078211
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_85
timestamp 1562078211
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_97
timestamp 1562078211
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_113
timestamp 1562078211
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_125
timestamp 1562078211
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_141
timestamp 1562078211
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_153
timestamp 1562078211
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_169
timestamp 1562078211
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_181
timestamp 1562078211
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_197
timestamp 1562078211
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_209
timestamp 1562078211
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_230
timestamp 1562078211
transform 1 0 22264 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_0_242
timestamp 1
transform 1 0 23368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_253
timestamp 1562078211
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_265
timestamp 1562078211
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_281
timestamp 1562078211
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_0_293
timestamp 1
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_3
timestamp 1562078211
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_15
timestamp 1562078211
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_27
timestamp 1562078211
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_39
timestamp 1562078211
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_57
timestamp 1562078211
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_69
timestamp 1562078211
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_81
timestamp 1562078211
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_93
timestamp 1562078211
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_109
timestamp 1
transform 1 0 11132 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_113
timestamp 1562078211
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_125
timestamp 1562078211
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_137
timestamp 1562078211
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_149
timestamp 1562078211
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_165
timestamp 1
transform 1 0 16284 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_169
timestamp 1562078211
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_181
timestamp 1562078211
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_193
timestamp 1562078211
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_205
timestamp 1562078211
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_225
timestamp 1562078211
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_237
timestamp 1562078211
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_249
timestamp 1562078211
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_261
timestamp 1562078211
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_277
timestamp 1
transform 1 0 26588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_281
timestamp 1562078211
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_293
timestamp 1
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 1
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_3
timestamp 1562078211
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_15
timestamp 1562078211
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_29
timestamp 1562078211
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_41
timestamp 1562078211
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_53
timestamp 1562078211
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_65
timestamp 1562078211
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 1
transform 1 0 8556 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_85
timestamp 1562078211
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_97
timestamp 1562078211
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_109
timestamp 1562078211
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_121
timestamp 1562078211
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_137
timestamp 1
transform 1 0 13708 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_141
timestamp 1562078211
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_153
timestamp 1562078211
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_165
timestamp 1562078211
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_177
timestamp 1562078211
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_193
timestamp 1
transform 1 0 18860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_197
timestamp 1562078211
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_209
timestamp 1562078211
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_221
timestamp 1562078211
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_233
timestamp 1562078211
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_249
timestamp 1
transform 1 0 24012 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_253
timestamp 1562078211
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_265
timestamp 1562078211
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_277
timestamp 1562078211
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_2_289
timestamp 1
transform 1 0 27692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_3
timestamp 1562078211
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_15
timestamp 1562078211
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_27
timestamp 1562078211
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_39
timestamp 1562078211
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_57
timestamp 1562078211
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_69
timestamp 1562078211
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_81
timestamp 1562078211
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_93
timestamp 1562078211
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1
transform 1 0 11132 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_113
timestamp 1562078211
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_125
timestamp 1562078211
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_137
timestamp 1562078211
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_149
timestamp 1562078211
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1
transform 1 0 16284 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_169
timestamp 1562078211
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_181
timestamp 1562078211
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_193
timestamp 1562078211
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_205
timestamp 1562078211
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_225
timestamp 1562078211
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_237
timestamp 1562078211
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_249
timestamp 1562078211
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_261
timestamp 1562078211
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_277
timestamp 1
transform 1 0 26588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_281
timestamp 1562078211
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_293
timestamp 1
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_297
timestamp 1
transform 1 0 28428 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_3
timestamp 1562078211
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_15
timestamp 1562078211
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_29
timestamp 1562078211
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_41
timestamp 1562078211
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_53
timestamp 1562078211
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_65
timestamp 1562078211
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1
transform 1 0 8556 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_85
timestamp 1562078211
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_97
timestamp 1562078211
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_109
timestamp 1562078211
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_121
timestamp 1562078211
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1
transform 1 0 13708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_141
timestamp 1562078211
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_153
timestamp 1562078211
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_165
timestamp 1562078211
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_177
timestamp 1562078211
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1
transform 1 0 18860 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_197
timestamp 1562078211
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_209
timestamp 1562078211
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_221
timestamp 1562078211
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_233
timestamp 1562078211
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_249
timestamp 1
transform 1 0 24012 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_253
timestamp 1562078211
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_265
timestamp 1562078211
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_277
timestamp 1562078211
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_4_289
timestamp 1
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_3
timestamp 1562078211
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_15
timestamp 1562078211
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_27
timestamp 1562078211
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_39
timestamp 1562078211
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_57
timestamp 1562078211
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_69
timestamp 1562078211
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_81
timestamp 1562078211
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_93
timestamp 1562078211
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1
transform 1 0 11132 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_113
timestamp 1562078211
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_125
timestamp 1562078211
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_137
timestamp 1562078211
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_149
timestamp 1562078211
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1
transform 1 0 16284 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_169
timestamp 1562078211
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_181
timestamp 1562078211
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_193
timestamp 1562078211
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_205
timestamp 1562078211
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1
transform 1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_225
timestamp 1562078211
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_237
timestamp 1562078211
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_249
timestamp 1562078211
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_261
timestamp 1562078211
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_277
timestamp 1
transform 1 0 26588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_281
timestamp 1562078211
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_293
timestamp 1
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_3
timestamp 1562078211
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_15
timestamp 1562078211
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_29
timestamp 1562078211
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_41
timestamp 1562078211
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_53
timestamp 1562078211
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_65
timestamp 1562078211
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_81
timestamp 1
transform 1 0 8556 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_85
timestamp 1562078211
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_97
timestamp 1562078211
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_109
timestamp 1562078211
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_121
timestamp 1562078211
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_137
timestamp 1
transform 1 0 13708 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_141
timestamp 1562078211
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_153
timestamp 1562078211
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_165
timestamp 1562078211
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_177
timestamp 1562078211
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_193
timestamp 1
transform 1 0 18860 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_197
timestamp 1562078211
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_209
timestamp 1562078211
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_221
timestamp 1562078211
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_233
timestamp 1562078211
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_249
timestamp 1
transform 1 0 24012 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_253
timestamp 1562078211
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_265
timestamp 1562078211
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_277
timestamp 1562078211
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_6_289
timestamp 1
transform 1 0 27692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_3
timestamp 1562078211
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_15
timestamp 1562078211
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_27
timestamp 1562078211
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_39
timestamp 1562078211
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_57
timestamp 1562078211
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_69
timestamp 1562078211
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_81
timestamp 1562078211
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_93
timestamp 1562078211
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1
transform 1 0 11132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_113
timestamp 1562078211
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_125
timestamp 1562078211
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_137
timestamp 1562078211
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_149
timestamp 1562078211
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_165
timestamp 1
transform 1 0 16284 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_169
timestamp 1562078211
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_181
timestamp 1562078211
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_193
timestamp 1562078211
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_205
timestamp 1562078211
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_225
timestamp 1562078211
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_237
timestamp 1562078211
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_249
timestamp 1562078211
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_261
timestamp 1562078211
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_277
timestamp 1
transform 1 0 26588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_281
timestamp 1562078211
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_293
timestamp 1
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 1
transform 1 0 28428 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_3
timestamp 1562078211
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_15
timestamp 1562078211
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_29
timestamp 1562078211
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_41
timestamp 1562078211
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_53
timestamp 1562078211
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_65
timestamp 1562078211
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_81
timestamp 1
transform 1 0 8556 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_85
timestamp 1562078211
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_97
timestamp 1562078211
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_109
timestamp 1562078211
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_121
timestamp 1562078211
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1
transform 1 0 13708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_141
timestamp 1562078211
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_153
timestamp 1562078211
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_165
timestamp 1562078211
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_177
timestamp 1562078211
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_193
timestamp 1
transform 1 0 18860 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_197
timestamp 1562078211
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_209
timestamp 1562078211
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_221
timestamp 1562078211
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_233
timestamp 1562078211
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_249
timestamp 1
transform 1 0 24012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_253
timestamp 1562078211
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_265
timestamp 1562078211
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_277
timestamp 1562078211
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_8_289
timestamp 1
transform 1 0 27692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_3
timestamp 1562078211
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_15
timestamp 1562078211
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_27
timestamp 1562078211
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_39
timestamp 1562078211
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_51
timestamp 1
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_57
timestamp 1562078211
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_69
timestamp 1562078211
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_81
timestamp 1562078211
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_93
timestamp 1562078211
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_105
timestamp 1
transform 1 0 10764 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1
transform 1 0 11132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_113
timestamp 1562078211
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_125
timestamp 1562078211
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_137
timestamp 1562078211
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_149
timestamp 1562078211
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_169
timestamp 1562078211
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_181
timestamp 1562078211
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_193
timestamp 1562078211
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_205
timestamp 1562078211
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_217
timestamp 1
transform 1 0 21068 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_225
timestamp 1562078211
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_237
timestamp 1562078211
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_249
timestamp 1562078211
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_261
timestamp 1562078211
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_273
timestamp 1
transform 1 0 26220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_277
timestamp 1
transform 1 0 26588 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_281
timestamp 1562078211
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_293
timestamp 1
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_297
timestamp 1
transform 1 0 28428 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_3
timestamp 1562078211
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_15
timestamp 1562078211
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_29
timestamp 1562078211
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_41
timestamp 1562078211
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_53
timestamp 1562078211
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_65
timestamp 1562078211
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_10_77
timestamp 1
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_81
timestamp 1
transform 1 0 8556 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_85
timestamp 1562078211
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_97
timestamp 1562078211
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_109
timestamp 1562078211
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_121
timestamp 1562078211
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_10_133
timestamp 1
transform 1 0 13340 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_137
timestamp 1
transform 1 0 13708 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_141
timestamp 1562078211
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_153
timestamp 1562078211
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_165
timestamp 1562078211
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_177
timestamp 1562078211
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_10_189
timestamp 1
transform 1 0 18492 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_193
timestamp 1
transform 1 0 18860 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_197
timestamp 1562078211
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_209
timestamp 1562078211
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_221
timestamp 1562078211
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_233
timestamp 1562078211
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_10_245
timestamp 1
transform 1 0 23644 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_249
timestamp 1
transform 1 0 24012 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_253
timestamp 1562078211
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_265
timestamp 1562078211
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_277
timestamp 1562078211
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_10_289
timestamp 1
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_293
timestamp 1
transform 1 0 28060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_295
timestamp 1
transform 1 0 28244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1
transform 1 0 28520 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_3
timestamp 1562078211
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_15
timestamp 1562078211
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_27
timestamp 1562078211
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_39
timestamp 1562078211
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_57
timestamp 1562078211
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_69
timestamp 1562078211
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_81
timestamp 1562078211
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_93
timestamp 1562078211
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_105
timestamp 1
transform 1 0 10764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1
transform 1 0 11132 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_113
timestamp 1562078211
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_125
timestamp 1562078211
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_137
timestamp 1562078211
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_149
timestamp 1562078211
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_161
timestamp 1
transform 1 0 15916 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_165
timestamp 1
transform 1 0 16284 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_169
timestamp 1562078211
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_181
timestamp 1562078211
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_193
timestamp 1562078211
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_205
timestamp 1562078211
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_217
timestamp 1
transform 1 0 21068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_225
timestamp 1562078211
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_237
timestamp 1562078211
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_249
timestamp 1562078211
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_261
timestamp 1562078211
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_273
timestamp 1
transform 1 0 26220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_277
timestamp 1
transform 1 0 26588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_281
timestamp 1
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_289
timestamp 1
transform 1 0 27692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_292
timestamp 1
transform 1 0 27968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_298
timestamp 1
transform 1 0 28520 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_3
timestamp 1562078211
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_15
timestamp 1562078211
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_29
timestamp 1562078211
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_41
timestamp 1562078211
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_53
timestamp 1562078211
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_65
timestamp 1562078211
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_77
timestamp 1
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_81
timestamp 1
transform 1 0 8556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_85
timestamp 1562078211
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_97
timestamp 1562078211
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_109
timestamp 1562078211
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_121
timestamp 1562078211
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_133
timestamp 1
transform 1 0 13340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_137
timestamp 1
transform 1 0 13708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_141
timestamp 1562078211
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_153
timestamp 1562078211
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_165
timestamp 1562078211
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_177
timestamp 1562078211
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_189
timestamp 1
transform 1 0 18492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1
transform 1 0 18860 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_197
timestamp 1562078211
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_209
timestamp 1562078211
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_221
timestamp 1562078211
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_233
timestamp 1562078211
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_245
timestamp 1
transform 1 0 23644 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_249
timestamp 1
transform 1 0 24012 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_253
timestamp 1562078211
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_265
timestamp 1562078211
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_277
timestamp 1562078211
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_12_289
timestamp 1
transform 1 0 27692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_3
timestamp 1562078211
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_15
timestamp 1562078211
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_27
timestamp 1562078211
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_39
timestamp 1562078211
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_57
timestamp 1562078211
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_69
timestamp 1562078211
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_81
timestamp 1562078211
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_93
timestamp 1562078211
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_105
timestamp 1
transform 1 0 10764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1
transform 1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_113
timestamp 1562078211
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_125
timestamp 1562078211
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_137
timestamp 1562078211
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_149
timestamp 1562078211
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_161
timestamp 1
transform 1 0 15916 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_13_164
timestamp 1
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_169
timestamp 1562078211
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_181
timestamp 1562078211
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_193
timestamp 1562078211
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_205
timestamp 1562078211
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_217
timestamp 1
transform 1 0 21068 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_225
timestamp 1562078211
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_237
timestamp 1562078211
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_249
timestamp 1562078211
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_261
timestamp 1562078211
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_273
timestamp 1
transform 1 0 26220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_277
timestamp 1
transform 1 0 26588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_281
timestamp 1562078211
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_293
timestamp 1
transform 1 0 28060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_3
timestamp 1562078211
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_15
timestamp 1562078211
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_29
timestamp 1562078211
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_41
timestamp 1562078211
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_53
timestamp 1562078211
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_65
timestamp 1562078211
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_14_77
timestamp 1
transform 1 0 8188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_81
timestamp 1
transform 1 0 8556 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_85
timestamp 1562078211
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_97
timestamp 1562078211
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_109
timestamp 1562078211
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_121
timestamp 1562078211
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_14_133
timestamp 1
transform 1 0 13340 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_137
timestamp 1
transform 1 0 13708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_141
timestamp 1562078211
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_14_153
timestamp 1
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_162
timestamp 1
transform 1 0 16008 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_180
timestamp 1562078211
transform 1 0 17664 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_14_192
timestamp 1
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_197
timestamp 1562078211
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_209
timestamp 1562078211
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_221
timestamp 1562078211
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_233
timestamp 1562078211
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_14_245
timestamp 1
transform 1 0 23644 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_249
timestamp 1
transform 1 0 24012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_253
timestamp 1562078211
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_265
timestamp 1562078211
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_277
timestamp 1562078211
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_14_289
timestamp 1
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_3
timestamp 1562078211
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_15
timestamp 1562078211
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_27
timestamp 1562078211
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_39
timestamp 1562078211
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_57
timestamp 1562078211
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_69
timestamp 1562078211
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_15_81
timestamp 1
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1
transform 1 0 9292 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_96
timestamp 1562078211
transform 1 0 9936 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_108
timestamp 1
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_113
timestamp 1562078211
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_15_125
timestamp 1
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_133
timestamp 1
transform 1 0 13340 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_152
timestamp 1562078211
transform 1 0 15088 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_164
timestamp 1
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_15_178
timestamp 1
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_190
timestamp 1562078211
transform 1 0 18584 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_202
timestamp 1
transform 1 0 19688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_204
timestamp 1
transform 1 0 19872 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_207
timestamp 1562078211
transform 1 0 20148 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_219
timestamp 1
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_225
timestamp 1562078211
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_237
timestamp 1562078211
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_249
timestamp 1562078211
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_261
timestamp 1562078211
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_273
timestamp 1
transform 1 0 26220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_277
timestamp 1
transform 1 0 26588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_281
timestamp 1562078211
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_293
timestamp 1
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_297
timestamp 1
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_3
timestamp 1562078211
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_15
timestamp 1562078211
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_29
timestamp 1562078211
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_16_41
timestamp 1
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp 1
transform 1 0 5244 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_16_63
timestamp 1
transform 1 0 6900 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_73
timestamp 1
transform 1 0 7820 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_79
timestamp 1
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_93
timestamp 1
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_104
timestamp 1562078211
transform 1 0 10672 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_16_116
timestamp 1
transform 1 0 11776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_122
timestamp 1
transform 1 0 12328 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_16_151
timestamp 1
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_171
timestamp 1
transform 1 0 16836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_182
timestamp 1
transform 1 0 17848 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_16_187
timestamp 1
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_197
timestamp 1
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_205
timestamp 1
transform 1 0 19964 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_16_215
timestamp 1
transform 1 0 20884 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_223
timestamp 1
transform 1 0 21620 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_229
timestamp 1
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_16_234
timestamp 1
transform 1 0 22632 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_238
timestamp 1
transform 1 0 23000 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_245
timestamp 1
transform 1 0 23644 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_249
timestamp 1
transform 1 0 24012 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_253
timestamp 1
transform 1 0 24380 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_256
timestamp 1562078211
transform 1 0 24656 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_268
timestamp 1562078211
transform 1 0 25760 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_280
timestamp 1562078211
transform 1 0 26864 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_16_292
timestamp 1
transform 1 0 27968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_296
timestamp 1
transform 1 0 28336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_298
timestamp 1
transform 1 0 28520 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_3
timestamp 1562078211
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_15
timestamp 1562078211
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_27
timestamp 1562078211
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_17_39
timestamp 1
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_52
timestamp 1
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_17_66
timestamp 1
transform 1 0 7176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_70
timestamp 1
transform 1 0 7544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_79
timestamp 1
transform 1 0 8372 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_17_97
timestamp 1
transform 1 0 10028 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_113
timestamp 1562078211
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_125
timestamp 1562078211
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_17_137
timestamp 1
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_141
timestamp 1
transform 1 0 14076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_148
timestamp 1
transform 1 0 14720 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_156
timestamp 1
transform 1 0 15456 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_165
timestamp 1
transform 1 0 16284 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_177
timestamp 1
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_185
timestamp 1562078211
transform 1 0 18124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_17_197
timestamp 1
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1
transform 1 0 21068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_233
timestamp 1
transform 1 0 22540 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_251
timestamp 1
transform 1 0 24196 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_253
timestamp 1
transform 1 0 24380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_259
timestamp 1
transform 1 0 24932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_268
timestamp 1562078211
transform 1 0 25760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_281
timestamp 1562078211
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_17_293
timestamp 1
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_3
timestamp 1562078211
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_15
timestamp 1562078211
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_29
timestamp 1562078211
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_18_41
timestamp 1
transform 1 0 4876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_65
timestamp 1
transform 1 0 7084 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_94
timestamp 1
transform 1 0 9752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_112
timestamp 1
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_18_130
timestamp 1
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_141
timestamp 1562078211
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_153
timestamp 1
transform 1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_155
timestamp 1
transform 1 0 15364 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1
transform 1 0 16100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_18_173
timestamp 1
transform 1 0 17020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_177
timestamp 1
transform 1 0 17388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_179
timestamp 1
transform 1 0 17572 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1
transform 1 0 20056 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_217
timestamp 1
transform 1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_227
timestamp 1
transform 1 0 21988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_237
timestamp 1
transform 1 0 22908 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_18_248
timestamp 1
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_253
timestamp 1
transform 1 0 24380 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_262
timestamp 1562078211
transform 1 0 25208 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_274
timestamp 1562078211
transform 1 0 26312 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_286
timestamp 1562078211
transform 1 0 27416 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_298
timestamp 1
transform 1 0 28520 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_3
timestamp 1562078211
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_15
timestamp 1562078211
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_27
timestamp 1562078211
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_19_39
timestamp 1
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp 1
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_49
timestamp 1
transform 1 0 5612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_59
timestamp 1
transform 1 0 6532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_65
timestamp 1
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_83
timestamp 1
transform 1 0 8740 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_19_93
timestamp 1
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_97
timestamp 1
transform 1 0 10028 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_19_107
timestamp 1
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_122
timestamp 1
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_130
timestamp 1562078211
transform 1 0 13064 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_142
timestamp 1562078211
transform 1 0 14168 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_19_154
timestamp 1
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1
transform 1 0 17572 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_187
timestamp 1
transform 1 0 18308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_19_192
timestamp 1
transform 1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_196
timestamp 1
transform 1 0 19136 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_204
timestamp 1
transform 1 0 19872 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_213
timestamp 1
transform 1 0 20700 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_225
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_19_232
timestamp 1
transform 1 0 22448 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_236
timestamp 1
transform 1 0 22816 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_244
timestamp 1
transform 1 0 23552 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_252
timestamp 1
transform 1 0 24288 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_260
timestamp 1562078211
transform 1 0 25024 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_19_272
timestamp 1
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_281
timestamp 1562078211
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_19_293
timestamp 1
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_3
timestamp 1562078211
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_15
timestamp 1562078211
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_29
timestamp 1562078211
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_41
timestamp 1562078211
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_20_53
timestamp 1
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_77
timestamp 1
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_81
timestamp 1
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_91
timestamp 1
transform 1 0 9476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_101
timestamp 1
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_119
timestamp 1562078211
transform 1 0 12052 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_20_131
timestamp 1
transform 1 0 13156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_144
timestamp 1562078211
transform 1 0 14352 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_20_156
timestamp 1
transform 1 0 15456 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_164
timestamp 1
transform 1 0 16192 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_172
timestamp 1
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_181
timestamp 1562078211
transform 1 0 17756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1
transform 1 0 18860 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_20_197
timestamp 1
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_209
timestamp 1
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_218
timestamp 1562078211
transform 1 0 21160 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_20_230
timestamp 1
transform 1 0 22264 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_245
timestamp 1
transform 1 0 23644 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_249
timestamp 1
transform 1 0 24012 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_253
timestamp 1562078211
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_265
timestamp 1562078211
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_277
timestamp 1562078211
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_20_289
timestamp 1
transform 1 0 27692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_3
timestamp 1562078211
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_15
timestamp 1562078211
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_27
timestamp 1562078211
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_39
timestamp 1562078211
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_21_51
timestamp 1
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_21_57
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_61
timestamp 1
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_21_71
timestamp 1
transform 1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_84
timestamp 1
transform 1 0 8832 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_101
timestamp 1
transform 1 0 10396 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_113
timestamp 1562078211
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_21_125
timestamp 1
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_145
timestamp 1
transform 1 0 14444 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_150
timestamp 1562078211
transform 1 0 14904 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_21_162
timestamp 1
transform 1 0 16008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_169
timestamp 1562078211
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_181
timestamp 1562078211
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_199
timestamp 1
transform 1 0 19412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_209
timestamp 1
transform 1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_21_219
timestamp 1
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_225
timestamp 1562078211
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_237
timestamp 1
transform 1 0 22908 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_239
timestamp 1
transform 1 0 23092 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_248
timestamp 1
transform 1 0 23920 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_257
timestamp 1562078211
transform 1 0 24748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_21_269
timestamp 1
transform 1 0 25852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_277
timestamp 1
transform 1 0 26588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_281
timestamp 1562078211
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_21_293
timestamp 1
transform 1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_3
timestamp 1562078211
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_15
timestamp 1562078211
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_29
timestamp 1562078211
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_41
timestamp 1562078211
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_53
timestamp 1562078211
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_22_65
timestamp 1
transform 1 0 7084 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1
transform 1 0 7452 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_75
timestamp 1
transform 1 0 8004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_22_85
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1
transform 1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_22_113
timestamp 1
transform 1 0 11500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_117
timestamp 1
transform 1 0 11868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_22_126
timestamp 1
transform 1 0 12696 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_137
timestamp 1
transform 1 0 13708 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_22_141
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_153
timestamp 1
transform 1 0 15180 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_158
timestamp 1562078211
transform 1 0 15640 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_170
timestamp 1562078211
transform 1 0 16744 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_182
timestamp 1562078211
transform 1 0 17848 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_197
timestamp 1
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_214
timestamp 1
transform 1 0 20792 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_22_224
timestamp 1
transform 1 0 21712 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_232
timestamp 1
transform 1 0 22448 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_234
timestamp 1
transform 1 0 22632 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_253
timestamp 1
transform 1 0 24380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_262
timestamp 1
transform 1 0 25208 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_267
timestamp 1562078211
transform 1 0 25668 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_279
timestamp 1562078211
transform 1 0 26772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_22_291
timestamp 1
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_298
timestamp 1
transform 1 0 28520 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_3
timestamp 1562078211
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_15
timestamp 1562078211
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_27
timestamp 1562078211
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_39
timestamp 1562078211
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_57
timestamp 1562078211
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_69
timestamp 1562078211
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_23_81
timestamp 1
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_95
timestamp 1562078211
transform 1 0 9844 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_107
timestamp 1
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_119
timestamp 1
transform 1 0 12052 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1
transform 1 0 13708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_155
timestamp 1562078211
transform 1 0 15364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_169
timestamp 1562078211
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_181
timestamp 1562078211
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_193
timestamp 1562078211
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_205
timestamp 1562078211
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_217
timestamp 1
transform 1 0 21068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_225
timestamp 1562078211
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_237
timestamp 1
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_241
timestamp 1
transform 1 0 23276 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_243
timestamp 1
transform 1 0 23460 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_247
timestamp 1
transform 1 0 23828 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_257
timestamp 1562078211
transform 1 0 24748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_23_269
timestamp 1
transform 1 0 25852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_277
timestamp 1
transform 1 0 26588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_281
timestamp 1562078211
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_293
timestamp 1
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1
transform 1 0 28428 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_3
timestamp 1562078211
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_15
timestamp 1562078211
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_29
timestamp 1562078211
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_41
timestamp 1562078211
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_53
timestamp 1562078211
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_65
timestamp 1562078211
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_24_77
timestamp 1
transform 1 0 8188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_81
timestamp 1
transform 1 0 8556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_85
timestamp 1562078211
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_24_97
timestamp 1
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1
transform 1 0 10396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_103
timestamp 1
transform 1 0 10580 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_24_130
timestamp 1
transform 1 0 13064 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_160
timestamp 1562078211
transform 1 0 15824 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_172
timestamp 1562078211
transform 1 0 16928 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_184
timestamp 1562078211
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_197
timestamp 1562078211
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_209
timestamp 1562078211
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_221
timestamp 1562078211
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_233
timestamp 1562078211
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_24_245
timestamp 1
transform 1 0 23644 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_249
timestamp 1
transform 1 0 24012 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_253
timestamp 1562078211
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_265
timestamp 1562078211
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_277
timestamp 1562078211
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_24_289
timestamp 1
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_3
timestamp 1562078211
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_15
timestamp 1562078211
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_27
timestamp 1562078211
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_39
timestamp 1562078211
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_25_51
timestamp 1
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_57
timestamp 1562078211
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_69
timestamp 1562078211
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_81
timestamp 1562078211
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_93
timestamp 1562078211
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_25_105
timestamp 1
transform 1 0 10764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_109
timestamp 1
transform 1 0 11132 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_121
timestamp 1
transform 1 0 12236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_138
timestamp 1
transform 1 0 13800 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1
transform 1 0 14444 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_150
timestamp 1562078211
transform 1 0 14904 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_25_162
timestamp 1
transform 1 0 16008 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_169
timestamp 1562078211
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_181
timestamp 1562078211
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_193
timestamp 1562078211
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_205
timestamp 1562078211
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_25_217
timestamp 1
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_225
timestamp 1562078211
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_237
timestamp 1562078211
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_251
timestamp 1562078211
transform 1 0 24196 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_263
timestamp 1562078211
transform 1 0 25300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_25_275
timestamp 1
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_281
timestamp 1
transform 1 0 26956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp 1
transform 1 0 28520 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_3
timestamp 1562078211
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_15
timestamp 1562078211
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_29
timestamp 1562078211
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_41
timestamp 1562078211
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_53
timestamp 1
transform 1 0 5980 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_77
timestamp 1
transform 1 0 8188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_81
timestamp 1
transform 1 0 8556 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_85
timestamp 1562078211
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_97
timestamp 1562078211
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_26_109
timestamp 1
transform 1 0 11132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_113
timestamp 1
transform 1 0 11500 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1
transform 1 0 11684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1
transform 1 0 12880 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_26_135
timestamp 1
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_141
timestamp 1562078211
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_153
timestamp 1562078211
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_165
timestamp 1562078211
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_177
timestamp 1562078211
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_26_189
timestamp 1
transform 1 0 18492 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_193
timestamp 1
transform 1 0 18860 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_197
timestamp 1562078211
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_209
timestamp 1562078211
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_221
timestamp 1562078211
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_26_233
timestamp 1
transform 1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_241
timestamp 1
transform 1 0 23276 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_249
timestamp 1
transform 1 0 24012 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_255
timestamp 1
transform 1 0 24564 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_272
timestamp 1562078211
transform 1 0 26128 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_284
timestamp 1
transform 1 0 27232 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_286
timestamp 1
transform 1 0 27416 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_290
timestamp 1
transform 1 0 27784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_26_294
timestamp 1
transform 1 0 28152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_298
timestamp 1
transform 1 0 28520 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1
transform 1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_11
timestamp 1562078211
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_23
timestamp 1
transform 1 0 3220 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_40
timestamp 1
transform 1 0 4784 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_42
timestamp 1
transform 1 0 4968 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_48
timestamp 1
transform 1 0 5520 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_27_57
timestamp 1
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_69
timestamp 1
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1
transform 1 0 7820 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_75
timestamp 1
transform 1 0 8004 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_92
timestamp 1
transform 1 0 9568 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_27_113
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_124
timestamp 1562078211
transform 1 0 12512 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_136
timestamp 1562078211
transform 1 0 13616 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_27_148
timestamp 1
transform 1 0 14720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_161
timestamp 1
transform 1 0 15916 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_165
timestamp 1
transform 1 0 16284 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_27_169
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_180
timestamp 1
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_186
timestamp 1
transform 1 0 18216 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1
transform 1 0 20240 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_27_215
timestamp 1
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_27_225
timestamp 1
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_234
timestamp 1
transform 1 0 22632 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_27_243
timestamp 1
transform 1 0 23460 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_251
timestamp 1
transform 1 0 24196 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_260
timestamp 1562078211
transform 1 0 25024 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_27_272
timestamp 1
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_281
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_3
timestamp 1562078211
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_28_15
timestamp 1
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_19
timestamp 1
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_25
timestamp 1
transform 1 0 3404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_29
timestamp 1
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_37
timestamp 1
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_54
timestamp 1
transform 1 0 6072 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_78
timestamp 1
transform 1 0 8280 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_28_85
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_94
timestamp 1
transform 1 0 9752 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp 1
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_118
timestamp 1
transform 1 0 11960 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_122
timestamp 1562078211
transform 1 0 12328 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_28_134
timestamp 1
transform 1 0 13432 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_28_141
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_158
timestamp 1
transform 1 0 15640 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_160
timestamp 1
transform 1 0 15824 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_28_178
timestamp 1
transform 1 0 17480 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_28_190
timestamp 1
transform 1 0 18584 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_204
timestamp 1
transform 1 0 19872 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_206
timestamp 1
transform 1 0 20056 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_214
timestamp 1
transform 1 0 20792 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_219
timestamp 1
transform 1 0 21252 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_221
timestamp 1
transform 1 0 21436 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_231
timestamp 1
transform 1 0 22356 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_239
timestamp 1
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_249
timestamp 1
transform 1 0 24012 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_253
timestamp 1
transform 1 0 24380 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_260
timestamp 1562078211
transform 1 0 25024 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_272
timestamp 1562078211
transform 1 0 26128 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_284
timestamp 1562078211
transform 1 0 27232 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_296
timestamp 1
transform 1 0 28336 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_298
timestamp 1
transform 1 0 28520 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_7
timestamp 1562078211
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_29_19
timestamp 1
transform 1 0 2852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp 1
transform 1 0 3588 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_37
timestamp 1
transform 1 0 4508 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_64
timestamp 1
transform 1 0 6992 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_74
timestamp 1
transform 1 0 7912 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_96
timestamp 1
transform 1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp 1
transform 1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_122
timestamp 1562078211
transform 1 0 12328 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_134
timestamp 1562078211
transform 1 0 13432 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_29_146
timestamp 1
transform 1 0 14536 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_154
timestamp 1
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1
transform 1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_169
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_178
timestamp 1
transform 1 0 17480 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_186
timestamp 1
transform 1 0 18216 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1
transform 1 0 20608 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_29_220
timestamp 1
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_225
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_232
timestamp 1
transform 1 0 22448 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_250
timestamp 1562078211
transform 1 0 24104 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_262
timestamp 1562078211
transform 1 0 25208 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_29_274
timestamp 1
transform 1 0 26312 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_281
timestamp 1562078211
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_29_293
timestamp 1
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_297
timestamp 1
transform 1 0 28428 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_3
timestamp 1562078211
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_15
timestamp 1562078211
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_31
timestamp 1
transform 1 0 3956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_37
timestamp 1
transform 1 0 4508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_61
timestamp 1
transform 1 0 6716 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_70
timestamp 1
transform 1 0 7544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_103
timestamp 1
transform 1 0 10580 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_113
timestamp 1562078211
transform 1 0 11500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_125
timestamp 1562078211
transform 1 0 12604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_137
timestamp 1
transform 1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_141
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_159
timestamp 1
transform 1 0 15732 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_177
timestamp 1
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 1
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_30_204
timestamp 1
transform 1 0 19872 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_208
timestamp 1
transform 1 0 20240 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_225
timestamp 1
transform 1 0 21804 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_243
timestamp 1
transform 1 0 23460 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_249
timestamp 1
transform 1 0 24012 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_253
timestamp 1
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_262
timestamp 1562078211
transform 1 0 25208 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_274
timestamp 1562078211
transform 1 0 26312 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_286
timestamp 1562078211
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_298
timestamp 1
transform 1 0 28520 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_3
timestamp 1562078211
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_15
timestamp 1562078211
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_27
timestamp 1562078211
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_31_39
timestamp 1
transform 1 0 4692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_52
timestamp 1
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_31_66
timestamp 1
transform 1 0 7176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1
transform 1 0 7544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_72
timestamp 1
transform 1 0 7728 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_89
timestamp 1
transform 1 0 9292 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_99
timestamp 1
transform 1 0 10212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_31_106
timestamp 1
transform 1 0 10856 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_113
timestamp 1562078211
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_31_125
timestamp 1
transform 1 0 12604 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_136
timestamp 1562078211
transform 1 0 13616 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_148
timestamp 1
transform 1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_150
timestamp 1
transform 1 0 14904 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_157
timestamp 1
transform 1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_31_163
timestamp 1
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp 1
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_31_178
timestamp 1
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_182
timestamp 1
transform 1 0 17848 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1
transform 1 0 18032 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_201
timestamp 1
transform 1 0 19596 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1
transform 1 0 20516 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_229
timestamp 1
transform 1 0 22172 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_239
timestamp 1
transform 1 0 23092 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_249
timestamp 1
transform 1 0 24012 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_253
timestamp 1562078211
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_265
timestamp 1562078211
transform 1 0 25484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_277
timestamp 1
transform 1 0 26588 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_281
timestamp 1562078211
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_31_293
timestamp 1
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1
transform 1 0 28428 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_3
timestamp 1562078211
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_15
timestamp 1562078211
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_29
timestamp 1562078211
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_32_41
timestamp 1
transform 1 0 4876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_51
timestamp 1
transform 1 0 5796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_58
timestamp 1
transform 1 0 6440 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_68
timestamp 1
transform 1 0 7360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_32_78
timestamp 1
transform 1 0 8280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_85
timestamp 1562078211
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_97
timestamp 1562078211
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_109
timestamp 1562078211
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_121
timestamp 1562078211
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_32_133
timestamp 1
transform 1 0 13340 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_137
timestamp 1
transform 1 0 13708 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_141
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_162
timestamp 1
transform 1 0 16008 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_32_168
timestamp 1
transform 1 0 16560 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_176
timestamp 1
transform 1 0 17296 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_183
timestamp 1
transform 1 0 17940 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_188
timestamp 1
transform 1 0 18400 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1
transform 1 0 19412 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_208
timestamp 1
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_212
timestamp 1
transform 1 0 20608 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_221
timestamp 1
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_233
timestamp 1
transform 1 0 22540 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_241
timestamp 1
transform 1 0 23276 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_32_245
timestamp 1
transform 1 0 23644 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_249
timestamp 1
transform 1 0 24012 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_253
timestamp 1562078211
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_265
timestamp 1562078211
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_277
timestamp 1562078211
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_32_289
timestamp 1
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_3
timestamp 1562078211
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_15
timestamp 1562078211
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_27
timestamp 1562078211
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_39
timestamp 1562078211
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_33_51
timestamp 1
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_74
timestamp 1562078211
transform 1 0 7912 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_86
timestamp 1562078211
transform 1 0 9016 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_98
timestamp 1562078211
transform 1 0 10120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_33_113
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1
transform 1 0 11868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_124
timestamp 1
transform 1 0 12512 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_128
timestamp 1562078211
transform 1 0 12880 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_33_140
timestamp 1
transform 1 0 13984 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_144
timestamp 1
transform 1 0 14352 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_33_162
timestamp 1
transform 1 0 16008 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_169
timestamp 1562078211
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_181
timestamp 1562078211
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_33_193
timestamp 1
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1
transform 1 0 19596 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_33_208
timestamp 1
transform 1 0 20240 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_216
timestamp 1
transform 1 0 20976 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_225
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_231
timestamp 1
transform 1 0 22356 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_236
timestamp 1562078211
transform 1 0 22816 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_248
timestamp 1562078211
transform 1 0 23920 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_260
timestamp 1562078211
transform 1 0 25024 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_33_272
timestamp 1
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_281
timestamp 1562078211
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_33_293
timestamp 1
transform 1 0 28060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1
transform 1 0 28428 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_3
timestamp 1562078211
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_15
timestamp 1562078211
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_29
timestamp 1562078211
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_41
timestamp 1562078211
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_53
timestamp 1562078211
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_65
timestamp 1562078211
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_34_77
timestamp 1
transform 1 0 8188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_81
timestamp 1
transform 1 0 8556 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_85
timestamp 1562078211
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_34_97
timestamp 1
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_101
timestamp 1
transform 1 0 10396 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_118
timestamp 1
transform 1 0 11960 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_34_136
timestamp 1
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_34_141
timestamp 1
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_149
timestamp 1
transform 1 0 14812 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_34_153
timestamp 1
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_165
timestamp 1562078211
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_177
timestamp 1562078211
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_34_189
timestamp 1
transform 1 0 18492 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_193
timestamp 1
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_197
timestamp 1562078211
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_209
timestamp 1562078211
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_221
timestamp 1562078211
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_233
timestamp 1562078211
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_34_245
timestamp 1
transform 1 0 23644 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_249
timestamp 1
transform 1 0 24012 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_253
timestamp 1562078211
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_265
timestamp 1562078211
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_277
timestamp 1562078211
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_34_289
timestamp 1
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_3
timestamp 1562078211
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_15
timestamp 1562078211
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_27
timestamp 1562078211
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_39
timestamp 1562078211
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_51
timestamp 1
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_57
timestamp 1562078211
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_69
timestamp 1562078211
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_81
timestamp 1562078211
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_93
timestamp 1
transform 1 0 9660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_97
timestamp 1
transform 1 0 10028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_99
timestamp 1
transform 1 0 10212 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_102
timestamp 1
transform 1 0 10488 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_109
timestamp 1
transform 1 0 11132 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp 1
transform 1 0 12144 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1
transform 1 0 12880 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_132
timestamp 1562078211
transform 1 0 13248 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_144
timestamp 1562078211
transform 1 0 14352 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_156
timestamp 1562078211
transform 1 0 15456 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_169
timestamp 1562078211
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_181
timestamp 1562078211
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_193
timestamp 1562078211
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_205
timestamp 1562078211
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_217
timestamp 1
transform 1 0 21068 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_221
timestamp 1
transform 1 0 21436 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_225
timestamp 1562078211
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_237
timestamp 1562078211
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_249
timestamp 1562078211
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_261
timestamp 1562078211
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_273
timestamp 1
transform 1 0 26220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_277
timestamp 1
transform 1 0 26588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_281
timestamp 1562078211
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_293
timestamp 1
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_297
timestamp 1
transform 1 0 28428 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_3
timestamp 1
transform 1 0 1380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_7
timestamp 1
transform 1 0 1748 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_11
timestamp 1562078211
transform 1 0 2116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_36_23
timestamp 1
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_29
timestamp 1562078211
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_41
timestamp 1562078211
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_53
timestamp 1562078211
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_65
timestamp 1562078211
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_36_77
timestamp 1
transform 1 0 8188 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_81
timestamp 1
transform 1 0 8556 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_85
timestamp 1
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_93
timestamp 1
transform 1 0 9660 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1
transform 1 0 10488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_36_109
timestamp 1
transform 1 0 11132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_121
timestamp 1
transform 1 0 12236 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_150
timestamp 1562078211
transform 1 0 14904 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_36_162
timestamp 1
transform 1 0 16008 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_170
timestamp 1
transform 1 0 16744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_173
timestamp 1
transform 1 0 17020 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_197
timestamp 1562078211
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_209
timestamp 1562078211
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_221
timestamp 1562078211
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_36_233
timestamp 1
transform 1 0 22540 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_237
timestamp 1
transform 1 0 22908 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_36_242
timestamp 1
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_253
timestamp 1562078211
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_265
timestamp 1562078211
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_277
timestamp 1562078211
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_36_289
timestamp 1
transform 1 0 27692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_3
timestamp 1562078211
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_15
timestamp 1562078211
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_37_27
timestamp 1
transform 1 0 3588 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_31
timestamp 1
transform 1 0 3956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_33
timestamp 1
transform 1 0 4140 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_39
timestamp 1
transform 1 0 4692 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_43
timestamp 1562078211
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_57
timestamp 1562078211
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_37_69
timestamp 1
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_77
timestamp 1
transform 1 0 8188 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_83
timestamp 1
transform 1 0 8740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_87
timestamp 1
transform 1 0 9108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_89
timestamp 1
transform 1 0 9292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_106
timestamp 1
transform 1 0 10856 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_108
timestamp 1
transform 1 0 11040 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_122
timestamp 1
transform 1 0 12328 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_124
timestamp 1
transform 1 0 12512 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_141
timestamp 1
transform 1 0 14076 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_151
timestamp 1562078211
transform 1 0 14996 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_37_163
timestamp 1
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_169
timestamp 1562078211
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_37_181
timestamp 1
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_185
timestamp 1
transform 1 0 18124 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_190
timestamp 1
transform 1 0 18584 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_192
timestamp 1
transform 1 0 18768 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_201
timestamp 1
transform 1 0 19596 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_208
timestamp 1562078211
transform 1 0 20240 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_37_220
timestamp 1
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_225
timestamp 1
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_229
timestamp 1
transform 1 0 22172 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_247
timestamp 1
transform 1 0 23828 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_252
timestamp 1562078211
transform 1 0 24288 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_264
timestamp 1562078211
transform 1 0 25392 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_37_276
timestamp 1
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_281
timestamp 1562078211
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_37_293
timestamp 1
transform 1 0 28060 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_297
timestamp 1
transform 1 0 28428 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_3
timestamp 1562078211
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_15
timestamp 1562078211
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_29
timestamp 1562078211
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_38_41
timestamp 1
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_65
timestamp 1
transform 1 0 7084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_69
timestamp 1
transform 1 0 7452 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_71
timestamp 1
transform 1 0 7636 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_38_80
timestamp 1
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_87
timestamp 1
transform 1 0 9108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_104
timestamp 1
transform 1 0 10672 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_119
timestamp 1
transform 1 0 12052 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_130
timestamp 1
transform 1 0 13064 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_148
timestamp 1
transform 1 0 14720 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_38_152
timestamp 1
transform 1 0 15088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_156
timestamp 1
transform 1 0 15456 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_38_173
timestamp 1
transform 1 0 17020 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_177
timestamp 1
transform 1 0 17388 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_179
timestamp 1
transform 1 0 17572 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_184
timestamp 1
transform 1 0 18032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_197
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_214
timestamp 1
transform 1 0 20792 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1
transform 1 0 21252 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_38_237
timestamp 1
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_241
timestamp 1
transform 1 0 23276 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_253
timestamp 1
transform 1 0 24380 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_260
timestamp 1562078211
transform 1 0 25024 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_272
timestamp 1562078211
transform 1 0 26128 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_284
timestamp 1562078211
transform 1 0 27232 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_296
timestamp 1
transform 1 0 28336 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_298
timestamp 1
transform 1 0 28520 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1
transform 1 0 1380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_7
timestamp 1562078211
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_19
timestamp 1562078211
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_31
timestamp 1562078211
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_43
timestamp 1562078211
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_57
timestamp 1562078211
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_69
timestamp 1562078211
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_81
timestamp 1
transform 1 0 8556 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_98
timestamp 1
transform 1 0 10120 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_105
timestamp 1
transform 1 0 10764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_109
timestamp 1
transform 1 0 11132 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_113
timestamp 1
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_117
timestamp 1
transform 1 0 11868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_39_127
timestamp 1
transform 1 0 12788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_131
timestamp 1
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_137
timestamp 1
transform 1 0 13708 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_141
timestamp 1562078211
transform 1 0 14076 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_39_153
timestamp 1
transform 1 0 15180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_157
timestamp 1
transform 1 0 15548 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_161
timestamp 1
transform 1 0 15916 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_169
timestamp 1
transform 1 0 16652 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_186
timestamp 1
transform 1 0 18216 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_204
timestamp 1
transform 1 0 19872 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_225
timestamp 1
transform 1 0 21804 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_234
timestamp 1
transform 1 0 22632 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_244
timestamp 1
transform 1 0 23552 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_246
timestamp 1
transform 1 0 23736 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_263
timestamp 1562078211
transform 1 0 25300 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_39_275
timestamp 1
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_281
timestamp 1562078211
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_39_293
timestamp 1
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_297
timestamp 1
transform 1 0 28428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_7
timestamp 1562078211
transform 1 0 1748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_40_19
timestamp 1
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_29
timestamp 1562078211
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_41
timestamp 1562078211
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_53
timestamp 1562078211
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_65
timestamp 1562078211
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_40_77
timestamp 1
transform 1 0 8188 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_81
timestamp 1
transform 1 0 8556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_85
timestamp 1562078211
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_40_97
timestamp 1
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_40_109
timestamp 1
transform 1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_117
timestamp 1
transform 1 0 11868 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_126
timestamp 1562078211
transform 1 0 12696 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_141
timestamp 1562078211
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_153
timestamp 1562078211
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_165
timestamp 1
transform 1 0 16284 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_174
timestamp 1
transform 1 0 17112 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_40_182
timestamp 1
transform 1 0 17848 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_197
timestamp 1
transform 1 0 19228 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_40_206
timestamp 1
transform 1 0 20056 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_210
timestamp 1
transform 1 0 20424 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_219
timestamp 1
transform 1 0 21252 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_40_229
timestamp 1
transform 1 0 22172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_233
timestamp 1
transform 1 0 22540 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_242
timestamp 1
transform 1 0 23368 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_249
timestamp 1
transform 1 0 24012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_253
timestamp 1
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_258
timestamp 1
transform 1 0 24840 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_262
timestamp 1562078211
transform 1 0 25208 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_274
timestamp 1562078211
transform 1 0 26312 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_286
timestamp 1562078211
transform 1 0 27416 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_298
timestamp 1
transform 1 0 28520 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_3
timestamp 1562078211
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_15
timestamp 1562078211
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_27
timestamp 1562078211
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_39
timestamp 1562078211
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_41_51
timestamp 1
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_57
timestamp 1562078211
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_69
timestamp 1562078211
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_81
timestamp 1562078211
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_93
timestamp 1562078211
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_41_105
timestamp 1
transform 1 0 10764 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_109
timestamp 1
transform 1 0 11132 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_41_113
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_117
timestamp 1
transform 1 0 11868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_119
timestamp 1
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_136
timestamp 1562078211
transform 1 0 13616 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_148
timestamp 1562078211
transform 1 0 14720 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_41_160
timestamp 1
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_169
timestamp 1562078211
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_181
timestamp 1
transform 1 0 17756 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_183
timestamp 1
transform 1 0 17940 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_189
timestamp 1
transform 1 0 18492 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_197
timestamp 1
transform 1 0 19228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_204
timestamp 1
transform 1 0 19872 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_206
timestamp 1
transform 1 0 20056 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_213
timestamp 1
transform 1 0 20700 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_225
timestamp 1
transform 1 0 21804 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_232
timestamp 1
transform 1 0 22448 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_240
timestamp 1
transform 1 0 23184 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_247
timestamp 1562078211
transform 1 0 23828 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_259
timestamp 1562078211
transform 1 0 24932 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_41_271
timestamp 1
transform 1 0 26036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_281
timestamp 1562078211
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_41_293
timestamp 1
transform 1 0 28060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_297
timestamp 1
transform 1 0 28428 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_3
timestamp 1562078211
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_15
timestamp 1562078211
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_29
timestamp 1562078211
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_41
timestamp 1562078211
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_53
timestamp 1562078211
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_65
timestamp 1562078211
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_42_77
timestamp 1
transform 1 0 8188 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_81
timestamp 1
transform 1 0 8556 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_85
timestamp 1562078211
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_97
timestamp 1562078211
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_109
timestamp 1562078211
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_121
timestamp 1562078211
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_42_133
timestamp 1
transform 1 0 13340 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_137
timestamp 1
transform 1 0 13708 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_141
timestamp 1562078211
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_153
timestamp 1562078211
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_165
timestamp 1562078211
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_177
timestamp 1562078211
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_42_189
timestamp 1
transform 1 0 18492 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_193
timestamp 1
transform 1 0 18860 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_42_197
timestamp 1
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_201
timestamp 1
transform 1 0 19596 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_42_206
timestamp 1
transform 1 0 20056 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_214
timestamp 1
transform 1 0 20792 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_220
timestamp 1562078211
transform 1 0 21344 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_232
timestamp 1562078211
transform 1 0 22448 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_42_244
timestamp 1
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_253
timestamp 1562078211
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_265
timestamp 1562078211
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_277
timestamp 1562078211
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_42_289
timestamp 1
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_3
timestamp 1562078211
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_15
timestamp 1562078211
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_27
timestamp 1562078211
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_39
timestamp 1562078211
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_43_51
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_57
timestamp 1562078211
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_69
timestamp 1562078211
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_83
timestamp 1
transform 1 0 8740 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_85
timestamp 1
transform 1 0 8924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_91
timestamp 1
transform 1 0 9476 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_95
timestamp 1562078211
transform 1 0 9844 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_43_107
timestamp 1
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_113
timestamp 1
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_121
timestamp 1
transform 1 0 12236 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_124
timestamp 1
transform 1 0 12512 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_131
timestamp 1
transform 1 0 13156 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_141
timestamp 1562078211
transform 1 0 14076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_153
timestamp 1562078211
transform 1 0 15180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_165
timestamp 1
transform 1 0 16284 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_169
timestamp 1562078211
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_43_181
timestamp 1
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_189
timestamp 1
transform 1 0 18492 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_191
timestamp 1
transform 1 0 18676 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_199
timestamp 1562078211
transform 1 0 19412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_211
timestamp 1562078211
transform 1 0 20516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_225
timestamp 1562078211
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_237
timestamp 1562078211
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_249
timestamp 1562078211
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_261
timestamp 1
transform 1 0 25116 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_270
timestamp 1
transform 1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_281
timestamp 1562078211
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_43_293
timestamp 1
transform 1 0 28060 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_297
timestamp 1
transform 1 0 28428 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_3
timestamp 1562078211
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_15
timestamp 1562078211
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_29
timestamp 1562078211
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_41
timestamp 1562078211
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_53
timestamp 1562078211
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_44_65
timestamp 1
transform 1 0 7084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_73
timestamp 1
transform 1 0 7820 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_75
timestamp 1
transform 1 0 8004 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_81
timestamp 1
transform 1 0 8556 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_85
timestamp 1
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_94
timestamp 1562078211
transform 1 0 9752 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_106
timestamp 1562078211
transform 1 0 10856 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_44_118
timestamp 1
transform 1 0 11960 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_122
timestamp 1
transform 1 0 12328 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_141
timestamp 1562078211
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_153
timestamp 1562078211
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_44_165
timestamp 1
transform 1 0 16284 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_173
timestamp 1
transform 1 0 17020 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_181
timestamp 1
transform 1 0 17756 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_44_190
timestamp 1
transform 1 0 18584 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_44_197
timestamp 1
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_201
timestamp 1
transform 1 0 19596 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_203
timestamp 1
transform 1 0 19780 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_213
timestamp 1562078211
transform 1 0 20700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_44_225
timestamp 1
transform 1 0 21804 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_229
timestamp 1
transform 1 0 22172 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_235
timestamp 1562078211
transform 1 0 22724 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_44_247
timestamp 1
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_253
timestamp 1562078211
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_265
timestamp 1562078211
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_277
timestamp 1562078211
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_44_289
timestamp 1
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_3
timestamp 1562078211
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_15
timestamp 1562078211
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_27
timestamp 1562078211
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_39
timestamp 1562078211
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_45_57
timestamp 1
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_61
timestamp 1
transform 1 0 6716 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_63
timestamp 1
transform 1 0 6900 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_80
timestamp 1
transform 1 0 8464 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_45_98
timestamp 1
transform 1 0 10120 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_109
timestamp 1
transform 1 0 11132 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_45_113
timestamp 1
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_117
timestamp 1
transform 1 0 11868 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_124
timestamp 1
transform 1 0 12512 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_45_128
timestamp 1
transform 1 0 12880 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_140
timestamp 1
transform 1 0 13984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_45_155
timestamp 1
transform 1 0 15364 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_163
timestamp 1
transform 1 0 16100 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_169
timestamp 1
transform 1 0 16652 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_178
timestamp 1
transform 1 0 17480 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_186
timestamp 1
transform 1 0 18216 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_193
timestamp 1562078211
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_205
timestamp 1562078211
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_45_217
timestamp 1
transform 1 0 21068 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_221
timestamp 1
transform 1 0 21436 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_225
timestamp 1
transform 1 0 21804 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_234
timestamp 1
transform 1 0 22632 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_243
timestamp 1
transform 1 0 23460 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_245
timestamp 1
transform 1 0 23644 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_255
timestamp 1
transform 1 0 24564 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_263
timestamp 1562078211
transform 1 0 25300 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_45_275
timestamp 1
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_281
timestamp 1562078211
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_45_293
timestamp 1
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1
transform 1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_3
timestamp 1562078211
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_15
timestamp 1562078211
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_29
timestamp 1562078211
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_41
timestamp 1562078211
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_46_53
timestamp 1
transform 1 0 5980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_57
timestamp 1
transform 1 0 6348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_74
timestamp 1
transform 1 0 7912 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_76
timestamp 1
transform 1 0 8096 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_85
timestamp 1
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_89
timestamp 1
transform 1 0 9292 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_98
timestamp 1
transform 1 0 10120 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_46_108
timestamp 1
transform 1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_112
timestamp 1
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_121
timestamp 1
transform 1 0 12236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_125
timestamp 1
transform 1 0 12604 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_134
timestamp 1
transform 1 0 13432 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_141
timestamp 1
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_144
timestamp 1
transform 1 0 14352 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_148
timestamp 1
transform 1 0 14720 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_165
timestamp 1
transform 1 0 16284 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_176
timestamp 1
transform 1 0 17296 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_183
timestamp 1
transform 1 0 17940 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_46_188
timestamp 1
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_197
timestamp 1562078211
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_46_209
timestamp 1
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_213
timestamp 1
transform 1 0 20700 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_230
timestamp 1
transform 1 0 22264 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_234
timestamp 1
transform 1 0 22632 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_253
timestamp 1
transform 1 0 24380 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_262
timestamp 1562078211
transform 1 0 25208 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_274
timestamp 1562078211
transform 1 0 26312 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_46_286
timestamp 1
transform 1 0 27416 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_294
timestamp 1
transform 1 0 28152 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_298
timestamp 1
transform 1 0 28520 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_3
timestamp 1562078211
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_15
timestamp 1562078211
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_27
timestamp 1562078211
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_39
timestamp 1562078211
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_57
timestamp 1
transform 1 0 6348 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_63
timestamp 1
transform 1 0 6900 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_65
timestamp 1
transform 1 0 7084 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_82
timestamp 1
transform 1 0 8648 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_47_92
timestamp 1
transform 1 0 9568 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_104
timestamp 1
transform 1 0 10672 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_113
timestamp 1
transform 1 0 11500 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_130
timestamp 1
transform 1 0 13064 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_139
timestamp 1
transform 1 0 13892 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_161
timestamp 1
transform 1 0 15916 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_165
timestamp 1
transform 1 0 16284 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_169
timestamp 1
transform 1 0 16652 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_179
timestamp 1
transform 1 0 17572 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_186
timestamp 1562078211
transform 1 0 18216 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_198
timestamp 1562078211
transform 1 0 19320 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_210
timestamp 1
transform 1 0 20424 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_213
timestamp 1
transform 1 0 20700 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_218
timestamp 1
transform 1 0 21160 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_227
timestamp 1
transform 1 0 21988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_47_236
timestamp 1
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_240
timestamp 1
transform 1 0 23184 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_244
timestamp 1
transform 1 0 23552 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_255
timestamp 1
transform 1 0 24564 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_260
timestamp 1
transform 1 0 25024 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_264
timestamp 1562078211
transform 1 0 25392 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_47_276
timestamp 1
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_281
timestamp 1562078211
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_47_293
timestamp 1
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_297
timestamp 1
transform 1 0 28428 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_3
timestamp 1562078211
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_15
timestamp 1562078211
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_29
timestamp 1
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_53
timestamp 1
transform 1 0 5980 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_55
timestamp 1
transform 1 0 6164 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_64
timestamp 1
transform 1 0 6992 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_68
timestamp 1
transform 1 0 7360 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_75
timestamp 1
transform 1 0 8004 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_85
timestamp 1
transform 1 0 8924 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1
transform 1 0 9660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_111
timestamp 1
transform 1 0 11316 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_48_115
timestamp 1
transform 1 0 11684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_135
timestamp 1
transform 1 0 13524 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_141
timestamp 1
transform 1 0 14076 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_48_154
timestamp 1
transform 1 0 15272 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_158
timestamp 1
transform 1 0 15640 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_160
timestamp 1
transform 1 0 15824 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_169
timestamp 1
transform 1 0 16652 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_177
timestamp 1
transform 1 0 17388 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_183
timestamp 1562078211
transform 1 0 17940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_197
timestamp 1
transform 1 0 19228 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_48_201
timestamp 1
transform 1 0 19596 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_205
timestamp 1
transform 1 0 19964 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_207
timestamp 1
transform 1 0 20148 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_216
timestamp 1
transform 1 0 20976 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_227
timestamp 1562078211
transform 1 0 21988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_239
timestamp 1
transform 1 0 23092 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_242
timestamp 1
transform 1 0 23368 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_253
timestamp 1
transform 1 0 24380 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_262
timestamp 1
transform 1 0 25208 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_272
timestamp 1562078211
transform 1 0 26128 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_284
timestamp 1562078211
transform 1 0 27232 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_296
timestamp 1
transform 1 0 28336 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_298
timestamp 1
transform 1 0 28520 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_3
timestamp 1562078211
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_15
timestamp 1562078211
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_32
timestamp 1
transform 1 0 4048 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_36
timestamp 1562078211
transform 1 0 4416 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_49_48
timestamp 1
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_57
timestamp 1562078211
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_69
timestamp 1
transform 1 0 7452 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_72
timestamp 1
transform 1 0 7728 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_79
timestamp 1
transform 1 0 8372 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_49_89
timestamp 1
transform 1 0 9292 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_93
timestamp 1
transform 1 0 9660 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_113
timestamp 1
transform 1 0 11500 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_122
timestamp 1
transform 1 0 12328 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_130
timestamp 1
transform 1 0 13064 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_134
timestamp 1
transform 1 0 13432 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_136
timestamp 1
transform 1 0 13616 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_140
timestamp 1
transform 1 0 13984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_49_147
timestamp 1
transform 1 0 14628 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_151
timestamp 1
transform 1 0 14996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_155
timestamp 1
transform 1 0 15364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_157
timestamp 1
transform 1 0 15548 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_165
timestamp 1
transform 1 0 16284 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_169
timestamp 1
transform 1 0 16652 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_173
timestamp 1562078211
transform 1 0 17020 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_185
timestamp 1
transform 1 0 18124 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_194
timestamp 1
transform 1 0 18952 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_204
timestamp 1562078211
transform 1 0 19872 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_49_216
timestamp 1
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_225
timestamp 1562078211
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_242
timestamp 1
transform 1 0 23368 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_251
timestamp 1
transform 1 0 24196 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_49_259
timestamp 1
transform 1 0 24932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_281
timestamp 1562078211
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_49_293
timestamp 1
transform 1 0 28060 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_297
timestamp 1
transform 1 0 28428 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_3
timestamp 1
transform 1 0 1380 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_7
timestamp 1562078211
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_50_19
timestamp 1
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_29
timestamp 1562078211
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_41
timestamp 1562078211
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_53
timestamp 1562078211
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_65
timestamp 1562078211
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_77
timestamp 1
transform 1 0 8188 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_85
timestamp 1
transform 1 0 8924 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_102
timestamp 1
transform 1 0 10488 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_112
timestamp 1562078211
transform 1 0 11408 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_124
timestamp 1562078211
transform 1 0 12512 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_50_136
timestamp 1
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_141
timestamp 1562078211
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_153
timestamp 1
transform 1 0 15180 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_157
timestamp 1562078211
transform 1 0 15548 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_50_169
timestamp 1
transform 1 0 16652 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_177
timestamp 1
transform 1 0 17388 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_197
timestamp 1
transform 1 0 19228 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_207
timestamp 1562078211
transform 1 0 20148 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_219
timestamp 1562078211
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_231
timestamp 1562078211
transform 1 0 22356 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_243
timestamp 1
transform 1 0 23460 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_245
timestamp 1
transform 1 0 23644 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_253
timestamp 1
transform 1 0 24380 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_256
timestamp 1562078211
transform 1 0 24656 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_268
timestamp 1562078211
transform 1 0 25760 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_280
timestamp 1562078211
transform 1 0 26864 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_50_292
timestamp 1
transform 1 0 27968 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_296
timestamp 1
transform 1 0 28336 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_298
timestamp 1
transform 1 0 28520 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_3
timestamp 1
transform 1 0 1380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_7
timestamp 1
transform 1 0 1748 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_11
timestamp 1562078211
transform 1 0 2116 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_23
timestamp 1562078211
transform 1 0 3220 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_35
timestamp 1562078211
transform 1 0 4324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_51_47
timestamp 1
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_57
timestamp 1562078211
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_69
timestamp 1562078211
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_81
timestamp 1
transform 1 0 8556 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_51_85
timestamp 1
transform 1 0 8924 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_89
timestamp 1
transform 1 0 9292 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_98
timestamp 1562078211
transform 1 0 10120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_113
timestamp 1562078211
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_125
timestamp 1562078211
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_137
timestamp 1562078211
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_149
timestamp 1562078211
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_51_161
timestamp 1
transform 1 0 15916 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_165
timestamp 1
transform 1 0 16284 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_169
timestamp 1
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_173
timestamp 1
transform 1 0 17020 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_175
timestamp 1
transform 1 0 17204 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_179
timestamp 1
transform 1 0 17572 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_184
timestamp 1
transform 1 0 18032 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_191
timestamp 1
transform 1 0 18676 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_201
timestamp 1562078211
transform 1 0 19596 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_51_213
timestamp 1
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_221
timestamp 1
transform 1 0 21436 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_225
timestamp 1562078211
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_51_237
timestamp 1
transform 1 0 22908 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_245
timestamp 1
transform 1 0 23644 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_252
timestamp 1562078211
transform 1 0 24288 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_264
timestamp 1562078211
transform 1 0 25392 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_51_276
timestamp 1
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_281
timestamp 1562078211
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_51_293
timestamp 1
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 1
transform 1 0 28428 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_3
timestamp 1562078211
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_15
timestamp 1562078211
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_29
timestamp 1562078211
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_52_41
timestamp 1
transform 1 0 4876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_45
timestamp 1
transform 1 0 5244 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_47
timestamp 1
transform 1 0 5428 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_64
timestamp 1
transform 1 0 6992 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_68
timestamp 1562078211
transform 1 0 7360 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_52_80
timestamp 1
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_85
timestamp 1562078211
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_97
timestamp 1562078211
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_109
timestamp 1562078211
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_121
timestamp 1562078211
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_52_133
timestamp 1
transform 1 0 13340 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_137
timestamp 1
transform 1 0 13708 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_141
timestamp 1562078211
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_153
timestamp 1562078211
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_165
timestamp 1562078211
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_177
timestamp 1
transform 1 0 17388 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_52_181
timestamp 1
transform 1 0 17756 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_189
timestamp 1
transform 1 0 18492 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_197
timestamp 1562078211
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_209
timestamp 1562078211
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_221
timestamp 1562078211
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_233
timestamp 1562078211
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_52_245
timestamp 1
transform 1 0 23644 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_249
timestamp 1
transform 1 0 24012 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_253
timestamp 1562078211
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_265
timestamp 1562078211
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_277
timestamp 1562078211
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_52_289
timestamp 1
transform 1 0 27692 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_297
timestamp 1
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_3
timestamp 1562078211
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_15
timestamp 1562078211
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_27
timestamp 1562078211
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_39
timestamp 1562078211
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_53_51
timestamp 1
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_57
timestamp 1
transform 1 0 6348 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_63
timestamp 1
transform 1 0 6900 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_65
timestamp 1
transform 1 0 7084 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_74
timestamp 1562078211
transform 1 0 7912 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_86
timestamp 1562078211
transform 1 0 9016 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_98
timestamp 1562078211
transform 1 0 10120 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_113
timestamp 1562078211
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_125
timestamp 1562078211
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_137
timestamp 1562078211
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_149
timestamp 1562078211
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_53_161
timestamp 1
transform 1 0 15916 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_165
timestamp 1
transform 1 0 16284 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_169
timestamp 1562078211
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_181
timestamp 1562078211
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_193
timestamp 1562078211
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_53_205
timestamp 1
transform 1 0 19964 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_213
timestamp 1
transform 1 0 20700 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_215
timestamp 1
transform 1 0 20884 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_225
timestamp 1
transform 1 0 21804 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_231
timestamp 1562078211
transform 1 0 22356 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_243
timestamp 1562078211
transform 1 0 23460 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_255
timestamp 1562078211
transform 1 0 24564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_267
timestamp 1562078211
transform 1 0 25668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_281
timestamp 1562078211
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_53_293
timestamp 1
transform 1 0 28060 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 1
transform 1 0 28428 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_3
timestamp 1562078211
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_15
timestamp 1562078211
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_29
timestamp 1562078211
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_54_41
timestamp 1
transform 1 0 4876 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_45
timestamp 1
transform 1 0 5244 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_62
timestamp 1
transform 1 0 6808 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_72
timestamp 1
transform 1 0 7728 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_79
timestamp 1
transform 1 0 8372 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_85
timestamp 1562078211
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_97
timestamp 1562078211
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_109
timestamp 1562078211
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_54_121
timestamp 1
transform 1 0 12236 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_128
timestamp 1562078211
transform 1 0 12880 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_141
timestamp 1562078211
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_153
timestamp 1
transform 1 0 15180 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_163
timestamp 1
transform 1 0 16100 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_171
timestamp 1562078211
transform 1 0 16836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_54_183
timestamp 1
transform 1 0 17940 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_187
timestamp 1
transform 1 0 18308 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_189
timestamp 1
transform 1 0 18492 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_197
timestamp 1
transform 1 0 19228 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_54_205
timestamp 1
transform 1 0 19964 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_209
timestamp 1
transform 1 0 20332 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_214
timestamp 1
transform 1 0 20792 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_222
timestamp 1
transform 1 0 21528 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_231
timestamp 1
transform 1 0 22356 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_54_238
timestamp 1
transform 1 0 23000 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_246
timestamp 1
transform 1 0 23736 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_248
timestamp 1
transform 1 0 23920 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_253
timestamp 1562078211
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_265
timestamp 1562078211
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_277
timestamp 1562078211
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_54_289
timestamp 1
transform 1 0 27692 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_293
timestamp 1
transform 1 0 28060 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_298
timestamp 1
transform 1 0 28520 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_7
timestamp 1562078211
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_19
timestamp 1562078211
transform 1 0 2852 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_31
timestamp 1562078211
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_43
timestamp 1
transform 1 0 5060 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_46
timestamp 1
transform 1 0 5336 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_53
timestamp 1
transform 1 0 5980 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_57
timestamp 1
transform 1 0 6348 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_74
timestamp 1562078211
transform 1 0 7912 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_55_86
timestamp 1
transform 1 0 9016 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_94
timestamp 1
transform 1 0 9752 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_55_98
timestamp 1
transform 1 0 10120 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_102
timestamp 1
transform 1 0 10488 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_104
timestamp 1
transform 1 0 10672 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_55_119
timestamp 1
transform 1 0 12052 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_139
timestamp 1562078211
transform 1 0 13892 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_169
timestamp 1
transform 1 0 16652 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_178
timestamp 1562078211
transform 1 0 17480 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_190
timestamp 1
transform 1 0 18584 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_197
timestamp 1562078211
transform 1 0 19228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_209
timestamp 1562078211
transform 1 0 20332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_221
timestamp 1
transform 1 0 21436 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_225
timestamp 1
transform 1 0 21804 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_233
timestamp 1
transform 1 0 22540 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_241
timestamp 1
transform 1 0 23276 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_249
timestamp 1
transform 1 0 24012 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_258
timestamp 1
transform 1 0 24840 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_263
timestamp 1
transform 1 0 25300 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_268
timestamp 1562078211
transform 1 0 25760 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_281
timestamp 1
transform 1 0 26956 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_298
timestamp 1
transform 1 0 28520 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_3
timestamp 1562078211
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_15
timestamp 1562078211
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_29
timestamp 1562078211
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_56_41
timestamp 1
transform 1 0 4876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_45
timestamp 1
transform 1 0 5244 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_53
timestamp 1
transform 1 0 5980 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_63
timestamp 1
transform 1 0 6900 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_56_76
timestamp 1
transform 1 0 8096 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_85
timestamp 1
transform 1 0 8924 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_56_93
timestamp 1
transform 1 0 9660 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_97
timestamp 1
transform 1 0 10028 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_56_107
timestamp 1
transform 1 0 10948 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_111
timestamp 1
transform 1 0 11316 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_113
timestamp 1
transform 1 0 11500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_121
timestamp 1
transform 1 0 12236 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_141
timestamp 1
transform 1 0 14076 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_146
timestamp 1
transform 1 0 14536 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_56_150
timestamp 1
transform 1 0 14904 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_162
timestamp 1
transform 1 0 16008 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_166
timestamp 1562078211
transform 1 0 16376 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_184
timestamp 1
transform 1 0 18032 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_193
timestamp 1
transform 1 0 18860 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_197
timestamp 1
transform 1 0 19228 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_201
timestamp 1
transform 1 0 19596 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_56_206
timestamp 1
transform 1 0 20056 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_214
timestamp 1
transform 1 0 20792 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_222
timestamp 1
transform 1 0 21528 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_56_233
timestamp 1
transform 1 0 22540 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_237
timestamp 1
transform 1 0 22908 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_56_247
timestamp 1
transform 1 0 23828 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_253
timestamp 1
transform 1 0 24380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_262
timestamp 1
transform 1 0 25208 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_271
timestamp 1562078211
transform 1 0 26036 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_283
timestamp 1562078211
transform 1 0 27140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_56_295
timestamp 1
transform 1 0 28244 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_3
timestamp 1562078211
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_15
timestamp 1562078211
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_27
timestamp 1562078211
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_57_39
timestamp 1
transform 1 0 4692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_57
timestamp 1
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_85
timestamp 1
transform 1 0 8924 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_57_89
timestamp 1
transform 1 0 9292 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_101
timestamp 1
transform 1 0 10396 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_121
timestamp 1
transform 1 0 12236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_131
timestamp 1
transform 1 0 13156 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_141
timestamp 1
transform 1 0 14076 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_149
timestamp 1
transform 1 0 14812 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_169
timestamp 1562078211
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_197
timestamp 1
transform 1 0 19228 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_202
timestamp 1562078211
transform 1 0 19688 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_214
timestamp 1
transform 1 0 20792 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_218
timestamp 1
transform 1 0 21160 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_225
timestamp 1
transform 1 0 21804 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_242
timestamp 1
transform 1 0 23368 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_247
timestamp 1
transform 1 0 23828 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_249
timestamp 1
transform 1 0 24012 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_266
timestamp 1
transform 1 0 25576 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_57_276
timestamp 1
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_281
timestamp 1562078211
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_57_293
timestamp 1
transform 1 0 28060 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_297
timestamp 1
transform 1 0 28428 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_3
timestamp 1562078211
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_15
timestamp 1562078211
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_58_29
timestamp 1
transform 1 0 3772 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_33
timestamp 1
transform 1 0 4140 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_58_50
timestamp 1
transform 1 0 5704 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_54
timestamp 1
transform 1 0 6072 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_56
timestamp 1
transform 1 0 6256 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_65
timestamp 1
transform 1 0 7084 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_85
timestamp 1
transform 1 0 8924 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_102
timestamp 1
transform 1 0 10488 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_58_117
timestamp 1
transform 1 0 11868 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_129
timestamp 1
transform 1 0 12972 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_58_141
timestamp 1
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_148
timestamp 1
transform 1 0 14720 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_58_166
timestamp 1
transform 1 0 16376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_176
timestamp 1
transform 1 0 17296 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_184
timestamp 1
transform 1 0 18032 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_197
timestamp 1
transform 1 0 19228 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_206
timestamp 1562078211
transform 1 0 20056 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_58_218
timestamp 1
transform 1 0 21160 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_222
timestamp 1
transform 1 0 21528 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_231
timestamp 1562078211
transform 1 0 22356 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_58_243
timestamp 1
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_253
timestamp 1
transform 1 0 24380 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_262
timestamp 1562078211
transform 1 0 25208 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_274
timestamp 1562078211
transform 1 0 26312 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_286
timestamp 1562078211
transform 1 0 27416 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_298
timestamp 1
transform 1 0 28520 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_3
timestamp 1562078211
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_15
timestamp 1562078211
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_27
timestamp 1562078211
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_39
timestamp 1
transform 1 0 4692 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_46
timestamp 1
transform 1 0 5336 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_59_50
timestamp 1
transform 1 0 5704 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_57
timestamp 1
transform 1 0 6348 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_65
timestamp 1
transform 1 0 7084 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_59_75
timestamp 1
transform 1 0 8004 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_91
timestamp 1
transform 1 0 9476 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_100
timestamp 1
transform 1 0 10304 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_59_107
timestamp 1
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_59_113
timestamp 1
transform 1 0 11500 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_117
timestamp 1
transform 1 0 11868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_126
timestamp 1
transform 1 0 12696 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_128
timestamp 1
transform 1 0 12880 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_131
timestamp 1
transform 1 0 13156 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_139
timestamp 1
transform 1 0 13892 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_141
timestamp 1
transform 1 0 14076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_59_145
timestamp 1
transform 1 0 14444 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_155
timestamp 1
transform 1 0 15364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_165
timestamp 1
transform 1 0 16284 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_169
timestamp 1
transform 1 0 16652 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_190
timestamp 1
transform 1 0 18584 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_200
timestamp 1562078211
transform 1 0 19504 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_212
timestamp 1562078211
transform 1 0 20608 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_225
timestamp 1562078211
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_237
timestamp 1562078211
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_249
timestamp 1562078211
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_261
timestamp 1562078211
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_59_273
timestamp 1
transform 1 0 26220 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_277
timestamp 1
transform 1 0 26588 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_281
timestamp 1562078211
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_59_293
timestamp 1
transform 1 0 28060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_297
timestamp 1
transform 1 0 28428 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_3
timestamp 1562078211
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_15
timestamp 1562078211
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_29
timestamp 1562078211
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_47
timestamp 1
transform 1 0 5428 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_56
timestamp 1
transform 1 0 6256 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_66
timestamp 1562078211
transform 1 0 7176 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_60_78
timestamp 1
transform 1 0 8280 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_85
timestamp 1
transform 1 0 8924 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_91
timestamp 1
transform 1 0 9476 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_95
timestamp 1562078211
transform 1 0 9844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_60_107
timestamp 1
transform 1 0 10948 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_121
timestamp 1562078211
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_60_133
timestamp 1
transform 1 0 13340 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_137
timestamp 1
transform 1 0 13708 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_60_141
timestamp 1
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_145
timestamp 1
transform 1 0 14444 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_147
timestamp 1
transform 1 0 14628 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_150
timestamp 1562078211
transform 1 0 14904 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_170
timestamp 1
transform 1 0 16744 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_60_174
timestamp 1
transform 1 0 17112 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_182
timestamp 1
transform 1 0 17848 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_60_186
timestamp 1
transform 1 0 18216 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_197
timestamp 1562078211
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_209
timestamp 1562078211
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_221
timestamp 1562078211
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_233
timestamp 1562078211
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_60_245
timestamp 1
transform 1 0 23644 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_249
timestamp 1
transform 1 0 24012 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_253
timestamp 1562078211
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_265
timestamp 1562078211
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_277
timestamp 1562078211
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_60_289
timestamp 1
transform 1 0 27692 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_297
timestamp 1
transform 1 0 28428 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_3
timestamp 1562078211
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_15
timestamp 1562078211
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_27
timestamp 1
transform 1 0 3588 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_31
timestamp 1
transform 1 0 3956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_38
timestamp 1
transform 1 0 4600 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_45
timestamp 1
transform 1 0 5244 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_57
timestamp 1
transform 1 0 6348 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_74
timestamp 1562078211
transform 1 0 7912 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_86
timestamp 1562078211
transform 1 0 9016 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_98
timestamp 1562078211
transform 1 0 10120 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_113
timestamp 1562078211
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_125
timestamp 1562078211
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_137
timestamp 1562078211
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_149
timestamp 1562078211
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_161
timestamp 1
transform 1 0 15916 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_169
timestamp 1
transform 1 0 16652 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_172
timestamp 1562078211
transform 1 0 16928 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_184
timestamp 1562078211
transform 1 0 18032 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_196
timestamp 1562078211
transform 1 0 19136 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_208
timestamp 1562078211
transform 1 0 20240 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_61_220
timestamp 1
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_225
timestamp 1562078211
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_237
timestamp 1562078211
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_249
timestamp 1562078211
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_261
timestamp 1562078211
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_61_273
timestamp 1
transform 1 0 26220 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_277
timestamp 1
transform 1 0 26588 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_281
timestamp 1562078211
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_61_293
timestamp 1
transform 1 0 28060 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_297
timestamp 1
transform 1 0 28428 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_3
timestamp 1562078211
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_15
timestamp 1562078211
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_29
timestamp 1562078211
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_43
timestamp 1
transform 1 0 5060 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_61
timestamp 1
transform 1 0 6716 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_71
timestamp 1562078211
transform 1 0 7636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_85
timestamp 1562078211
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_97
timestamp 1562078211
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_109
timestamp 1562078211
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_121
timestamp 1562078211
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_62_133
timestamp 1
transform 1 0 13340 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_137
timestamp 1
transform 1 0 13708 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_141
timestamp 1562078211
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_153
timestamp 1562078211
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_165
timestamp 1562078211
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_177
timestamp 1562078211
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_62_189
timestamp 1
transform 1 0 18492 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_193
timestamp 1
transform 1 0 18860 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_197
timestamp 1562078211
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_209
timestamp 1562078211
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_221
timestamp 1562078211
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_233
timestamp 1562078211
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_62_245
timestamp 1
transform 1 0 23644 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_249
timestamp 1
transform 1 0 24012 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_253
timestamp 1562078211
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_265
timestamp 1562078211
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_277
timestamp 1562078211
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_62_289
timestamp 1
transform 1 0 27692 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_297
timestamp 1
transform 1 0 28428 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_3
timestamp 1562078211
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_15
timestamp 1562078211
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_27
timestamp 1562078211
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_63_39
timestamp 1
transform 1 0 4692 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_63_48
timestamp 1
transform 1 0 5520 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_57
timestamp 1
transform 1 0 6348 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_66
timestamp 1562078211
transform 1 0 7176 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_78
timestamp 1562078211
transform 1 0 8280 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_90
timestamp 1562078211
transform 1 0 9384 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_63_102
timestamp 1
transform 1 0 10488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_63_113
timestamp 1
transform 1 0 11500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_124
timestamp 1
transform 1 0 12512 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_126
timestamp 1
transform 1 0 12696 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_130
timestamp 1562078211
transform 1 0 13064 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_142
timestamp 1562078211
transform 1 0 14168 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_63_154
timestamp 1
transform 1 0 15272 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_162
timestamp 1
transform 1 0 16008 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_169
timestamp 1
transform 1 0 16652 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_175
timestamp 1562078211
transform 1 0 17204 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_187
timestamp 1562078211
transform 1 0 18308 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_199
timestamp 1562078211
transform 1 0 19412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_211
timestamp 1562078211
transform 1 0 20516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_225
timestamp 1562078211
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_237
timestamp 1562078211
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_249
timestamp 1562078211
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_261
timestamp 1562078211
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_63_273
timestamp 1
transform 1 0 26220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_277
timestamp 1
transform 1 0 26588 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_281
timestamp 1562078211
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_63_293
timestamp 1
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_297
timestamp 1
transform 1 0 28428 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_3
timestamp 1562078211
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_15
timestamp 1562078211
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_29
timestamp 1562078211
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_41
timestamp 1
transform 1 0 4876 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_58
timestamp 1
transform 1 0 6440 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_62
timestamp 1
transform 1 0 6808 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_69
timestamp 1562078211
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_81
timestamp 1
transform 1 0 8556 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_85
timestamp 1
transform 1 0 8924 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_88
timestamp 1562078211
transform 1 0 9200 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_64_100
timestamp 1
transform 1 0 10304 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_104
timestamp 1
transform 1 0 10672 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_112
timestamp 1
transform 1 0 11408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_122
timestamp 1
transform 1 0 12328 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_64_131
timestamp 1
transform 1 0 13156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_141
timestamp 1
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_152
timestamp 1
transform 1 0 15088 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_162
timestamp 1
transform 1 0 16008 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_180
timestamp 1
transform 1 0 17664 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_182
timestamp 1
transform 1 0 17848 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_189
timestamp 1
transform 1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_193
timestamp 1
transform 1 0 18860 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_197
timestamp 1562078211
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_209
timestamp 1562078211
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_221
timestamp 1562078211
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_233
timestamp 1562078211
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_64_245
timestamp 1
transform 1 0 23644 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_249
timestamp 1
transform 1 0 24012 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_253
timestamp 1562078211
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_265
timestamp 1562078211
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_277
timestamp 1562078211
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_64_289
timestamp 1
transform 1 0 27692 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_297
timestamp 1
transform 1 0 28428 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_3
timestamp 1562078211
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_20
timestamp 1
transform 1 0 2944 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_65_38
timestamp 1
transform 1 0 4600 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_50
timestamp 1
transform 1 0 5704 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_65_57
timestamp 1
transform 1 0 6348 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_61
timestamp 1
transform 1 0 6716 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_83
timestamp 1
transform 1 0 8740 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_65_101
timestamp 1
transform 1 0 10396 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_105
timestamp 1
transform 1 0 10764 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_113
timestamp 1
transform 1 0 11500 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_65_122
timestamp 1
transform 1 0 12328 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_126
timestamp 1
transform 1 0 12696 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_135
timestamp 1
transform 1 0 13524 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_139
timestamp 1
transform 1 0 13892 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_141
timestamp 1
transform 1 0 14076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_149
timestamp 1
transform 1 0 14812 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_65_159
timestamp 1
transform 1 0 15732 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_169
timestamp 1
transform 1 0 16652 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_178
timestamp 1
transform 1 0 17480 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_188
timestamp 1
transform 1 0 18400 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_198
timestamp 1
transform 1 0 19320 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_205
timestamp 1562078211
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_65_217
timestamp 1
transform 1 0 21068 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_221
timestamp 1
transform 1 0 21436 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_225
timestamp 1562078211
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_237
timestamp 1562078211
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_249
timestamp 1562078211
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_261
timestamp 1562078211
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_65_273
timestamp 1
transform 1 0 26220 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_277
timestamp 1
transform 1 0 26588 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_281
timestamp 1562078211
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_65_293
timestamp 1
transform 1 0 28060 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_297
timestamp 1
transform 1 0 28428 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_3
timestamp 1
transform 1 0 1380 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_7
timestamp 1
transform 1 0 1748 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_11
timestamp 1562078211
transform 1 0 2116 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_66_23
timestamp 1
transform 1 0 3220 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_29
timestamp 1562078211
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_41
timestamp 1562078211
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_53
timestamp 1562078211
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_65
timestamp 1562078211
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_66_77
timestamp 1
transform 1 0 8188 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_81
timestamp 1
transform 1 0 8556 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_85
timestamp 1
transform 1 0 8924 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_91
timestamp 1
transform 1 0 9476 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_66_95
timestamp 1
transform 1 0 9844 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_99
timestamp 1
transform 1 0 10212 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_106
timestamp 1
transform 1 0 10856 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_124
timestamp 1
transform 1 0 12512 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_126
timestamp 1
transform 1 0 12696 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_66_135
timestamp 1
transform 1 0 13524 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_141
timestamp 1
transform 1 0 14076 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_158
timestamp 1
transform 1 0 15640 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_66_163
timestamp 1
transform 1 0 16100 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_169
timestamp 1
transform 1 0 16652 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_171
timestamp 1
transform 1 0 16836 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_177
timestamp 1
transform 1 0 17388 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_197
timestamp 1
transform 1 0 19228 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_206
timestamp 1562078211
transform 1 0 20056 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_218
timestamp 1562078211
transform 1 0 21160 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_230
timestamp 1562078211
transform 1 0 22264 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_66_242
timestamp 1
transform 1 0 23368 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_253
timestamp 1562078211
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_265
timestamp 1562078211
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_277
timestamp 1562078211
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_66_289
timestamp 1
transform 1 0 27692 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_297
timestamp 1
transform 1 0 28428 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_3
timestamp 1562078211
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_15
timestamp 1562078211
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_27
timestamp 1562078211
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_39
timestamp 1562078211
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_67_51
timestamp 1
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_57
timestamp 1562078211
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_77
timestamp 1
transform 1 0 8188 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_95
timestamp 1
transform 1 0 9844 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_105
timestamp 1
transform 1 0 10764 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_113
timestamp 1
transform 1 0 11500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_129
timestamp 1
transform 1 0 12972 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_137
timestamp 1
transform 1 0 13708 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_142
timestamp 1
transform 1 0 14168 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_144
timestamp 1
transform 1 0 14352 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_153
timestamp 1
transform 1 0 15180 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_157
timestamp 1
transform 1 0 15548 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_164
timestamp 1
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_169
timestamp 1
transform 1 0 16652 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_177
timestamp 1
transform 1 0 17388 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_181
timestamp 1
transform 1 0 17756 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_198
timestamp 1
transform 1 0 19320 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_203
timestamp 1
transform 1 0 19780 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_208
timestamp 1
transform 1 0 20240 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_212
timestamp 1
transform 1 0 20608 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_67_216
timestamp 1
transform 1 0 20976 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_225
timestamp 1562078211
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_237
timestamp 1562078211
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_249
timestamp 1562078211
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_261
timestamp 1562078211
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_67_273
timestamp 1
transform 1 0 26220 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_277
timestamp 1
transform 1 0 26588 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_281
timestamp 1562078211
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_67_293
timestamp 1
transform 1 0 28060 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_297
timestamp 1
transform 1 0 28428 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_3
timestamp 1562078211
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_15
timestamp 1562078211
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_29
timestamp 1562078211
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_68_41
timestamp 1
transform 1 0 4876 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_65
timestamp 1
transform 1 0 7084 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_72
timestamp 1
transform 1 0 7728 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_74
timestamp 1
transform 1 0 7912 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_85
timestamp 1
transform 1 0 8924 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_91
timestamp 1
transform 1 0 9476 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_101
timestamp 1
transform 1 0 10396 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_68_110
timestamp 1
transform 1 0 11224 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_121
timestamp 1562078211
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_68_133
timestamp 1
transform 1 0 13340 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_137
timestamp 1
transform 1 0 13708 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_68_141
timestamp 1
transform 1 0 14076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_145
timestamp 1
transform 1 0 14444 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_153
timestamp 1
transform 1 0 15180 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_163
timestamp 1
transform 1 0 16100 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_165
timestamp 1
transform 1 0 16284 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_186
timestamp 1
transform 1 0 18216 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_197
timestamp 1
transform 1 0 19228 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_206
timestamp 1562078211
transform 1 0 20056 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_218
timestamp 1562078211
transform 1 0 21160 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_230
timestamp 1562078211
transform 1 0 22264 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_68_242
timestamp 1
transform 1 0 23368 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_253
timestamp 1562078211
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_265
timestamp 1562078211
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_277
timestamp 1562078211
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_68_289
timestamp 1
transform 1 0 27692 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_297
timestamp 1
transform 1 0 28428 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_3
timestamp 1562078211
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_15
timestamp 1562078211
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_27
timestamp 1562078211
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_39
timestamp 1562078211
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_69_51
timestamp 1
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_57
timestamp 1
transform 1 0 6348 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_61
timestamp 1
transform 1 0 6716 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_63
timestamp 1
transform 1 0 6900 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_72
timestamp 1
transform 1 0 7728 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_90
timestamp 1
transform 1 0 9384 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_69_108
timestamp 1
transform 1 0 11040 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_113
timestamp 1
transform 1 0 11500 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_121
timestamp 1562078211
transform 1 0 12236 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_69_133
timestamp 1
transform 1 0 13340 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_141
timestamp 1
transform 1 0 14076 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_69_148
timestamp 1
transform 1 0 14720 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_156
timestamp 1
transform 1 0 15456 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_163
timestamp 1
transform 1 0 16100 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_169
timestamp 1562078211
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_69_181
timestamp 1
transform 1 0 17756 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_185
timestamp 1
transform 1 0 18124 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_194
timestamp 1562078211
transform 1 0 18952 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_206
timestamp 1562078211
transform 1 0 20056 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_69_218
timestamp 1
transform 1 0 21160 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_225
timestamp 1562078211
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_237
timestamp 1562078211
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_249
timestamp 1562078211
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_261
timestamp 1562078211
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_69_273
timestamp 1
transform 1 0 26220 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_277
timestamp 1
transform 1 0 26588 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_281
timestamp 1562078211
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_69_293
timestamp 1
transform 1 0 28060 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_297
timestamp 1
transform 1 0 28428 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_3
timestamp 1562078211
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_15
timestamp 1562078211
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_29
timestamp 1562078211
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_70_41
timestamp 1
transform 1 0 4876 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_49
timestamp 1
transform 1 0 5612 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_51
timestamp 1
transform 1 0 5796 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_57
timestamp 1
transform 1 0 6348 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_59
timestamp 1
transform 1 0 6532 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_70_66
timestamp 1
transform 1 0 7176 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_70
timestamp 1
transform 1 0 7544 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_72
timestamp 1
transform 1 0 7728 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_70_79
timestamp 1
transform 1 0 8372 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_70_85
timestamp 1
transform 1 0 8924 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_89
timestamp 1
transform 1 0 9292 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_99
timestamp 1562078211
transform 1 0 10212 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_111
timestamp 1562078211
transform 1 0 11316 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_123
timestamp 1562078211
transform 1 0 12420 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_135
timestamp 1
transform 1 0 13524 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_141
timestamp 1562078211
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_153
timestamp 1
transform 1 0 15180 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_157
timestamp 1
transform 1 0 15548 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_159
timestamp 1
transform 1 0 15732 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_165
timestamp 1562078211
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_177
timestamp 1562078211
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_189
timestamp 1
transform 1 0 18492 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_193
timestamp 1
transform 1 0 18860 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_197
timestamp 1562078211
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_209
timestamp 1562078211
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_221
timestamp 1562078211
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_233
timestamp 1562078211
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_245
timestamp 1
transform 1 0 23644 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_249
timestamp 1
transform 1 0 24012 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_253
timestamp 1562078211
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_265
timestamp 1562078211
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_277
timestamp 1562078211
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_70_289
timestamp 1
transform 1 0 27692 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_297
timestamp 1
transform 1 0 28428 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_3
timestamp 1562078211
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_15
timestamp 1562078211
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_27
timestamp 1562078211
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_57
timestamp 1
transform 1 0 6348 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_66
timestamp 1
transform 1 0 7176 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_75
timestamp 1562078211
transform 1 0 8004 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_87
timestamp 1562078211
transform 1 0 9108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_99
timestamp 1562078211
transform 1 0 10212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_113
timestamp 1562078211
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_125
timestamp 1562078211
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_137
timestamp 1562078211
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_149
timestamp 1562078211
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_161
timestamp 1
transform 1 0 15916 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_165
timestamp 1
transform 1 0 16284 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_169
timestamp 1562078211
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_181
timestamp 1562078211
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_193
timestamp 1562078211
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_205
timestamp 1562078211
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_217
timestamp 1
transform 1 0 21068 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_221
timestamp 1
transform 1 0 21436 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_225
timestamp 1562078211
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_237
timestamp 1562078211
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_249
timestamp 1562078211
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_261
timestamp 1562078211
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_273
timestamp 1
transform 1 0 26220 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_277
timestamp 1
transform 1 0 26588 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_281
timestamp 1562078211
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_293
timestamp 1
transform 1 0 28060 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_297
timestamp 1
transform 1 0 28428 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_3
timestamp 1562078211
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_15
timestamp 1562078211
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_29
timestamp 1562078211
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_72_41
timestamp 1
transform 1 0 4876 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_54
timestamp 1562078211
transform 1 0 6072 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_66
timestamp 1562078211
transform 1 0 7176 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_72_78
timestamp 1
transform 1 0 8280 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_82
timestamp 1
transform 1 0 8648 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_85
timestamp 1562078211
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_97
timestamp 1562078211
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_109
timestamp 1562078211
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_121
timestamp 1562078211
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_133
timestamp 1
transform 1 0 13340 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_138
timestamp 1
transform 1 0 13800 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_141
timestamp 1562078211
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_153
timestamp 1562078211
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_165
timestamp 1562078211
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_177
timestamp 1562078211
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_72_189
timestamp 1
transform 1 0 18492 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_193
timestamp 1
transform 1 0 18860 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_197
timestamp 1562078211
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_209
timestamp 1562078211
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_221
timestamp 1562078211
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_233
timestamp 1562078211
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_72_245
timestamp 1
transform 1 0 23644 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_249
timestamp 1
transform 1 0 24012 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_253
timestamp 1562078211
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_265
timestamp 1562078211
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_277
timestamp 1562078211
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_72_289
timestamp 1
transform 1 0 27692 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_297
timestamp 1
transform 1 0 28428 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_3
timestamp 1562078211
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_15
timestamp 1562078211
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_27
timestamp 1562078211
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_73_39
timestamp 1
transform 1 0 4692 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_52
timestamp 1
transform 1 0 5888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_57
timestamp 1
transform 1 0 6348 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_66
timestamp 1562078211
transform 1 0 7176 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_78
timestamp 1562078211
transform 1 0 8280 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_90
timestamp 1562078211
transform 1 0 9384 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_73_102
timestamp 1
transform 1 0 10488 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_113
timestamp 1562078211
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_125
timestamp 1562078211
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_137
timestamp 1562078211
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_149
timestamp 1562078211
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_161
timestamp 1
transform 1 0 15916 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_165
timestamp 1
transform 1 0 16284 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_169
timestamp 1562078211
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_181
timestamp 1562078211
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_193
timestamp 1
transform 1 0 18860 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_197
timestamp 1
transform 1 0 19228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_201
timestamp 1
transform 1 0 19596 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_205
timestamp 1562078211
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_217
timestamp 1
transform 1 0 21068 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_221
timestamp 1
transform 1 0 21436 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_225
timestamp 1562078211
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_237
timestamp 1562078211
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_249
timestamp 1562078211
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_261
timestamp 1562078211
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_273
timestamp 1
transform 1 0 26220 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_277
timestamp 1
transform 1 0 26588 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_281
timestamp 1562078211
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_293
timestamp 1
transform 1 0 28060 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_297
timestamp 1
transform 1 0 28428 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_3
timestamp 1562078211
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_15
timestamp 1562078211
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_29
timestamp 1562078211
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_41
timestamp 1
transform 1 0 4876 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_59
timestamp 1562078211
transform 1 0 6532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_71
timestamp 1562078211
transform 1 0 7636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_85
timestamp 1562078211
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_74_97
timestamp 1
transform 1 0 10028 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_105
timestamp 1
transform 1 0 10764 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_112
timestamp 1
transform 1 0 11408 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_121
timestamp 1
transform 1 0 12236 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_126
timestamp 1562078211
transform 1 0 12696 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_138
timestamp 1
transform 1 0 13800 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_141
timestamp 1
transform 1 0 14076 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_145
timestamp 1
transform 1 0 14444 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_153
timestamp 1
transform 1 0 15180 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_74_157
timestamp 1
transform 1 0 15548 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_161
timestamp 1
transform 1 0 15916 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_170
timestamp 1562078211
transform 1 0 16744 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_182
timestamp 1
transform 1 0 17848 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_185
timestamp 1
transform 1 0 18124 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_187
timestamp 1
transform 1 0 18308 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_194
timestamp 1
transform 1 0 18952 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_197
timestamp 1
transform 1 0 19228 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_206
timestamp 1562078211
transform 1 0 20056 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_218
timestamp 1562078211
transform 1 0 21160 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_230
timestamp 1562078211
transform 1 0 22264 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_74_242
timestamp 1
transform 1 0 23368 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_253
timestamp 1562078211
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_265
timestamp 1562078211
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_277
timestamp 1562078211
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_74_289
timestamp 1
transform 1 0 27692 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_297
timestamp 1
transform 1 0 28428 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_3
timestamp 1562078211
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_15
timestamp 1562078211
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_27
timestamp 1562078211
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_39
timestamp 1562078211
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_51
timestamp 1
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_57
timestamp 1
transform 1 0 6348 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_66
timestamp 1562078211
transform 1 0 7176 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_78
timestamp 1562078211
transform 1 0 8280 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_75_90
timestamp 1
transform 1 0 9384 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_98
timestamp 1
transform 1 0 10120 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_100
timestamp 1
transform 1 0 10304 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_109
timestamp 1
transform 1 0 11132 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_113
timestamp 1
transform 1 0 11500 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_122
timestamp 1
transform 1 0 12328 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_75_127
timestamp 1
transform 1 0 12788 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_136
timestamp 1
transform 1 0 13616 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_75_145
timestamp 1
transform 1 0 14444 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_161
timestamp 1
transform 1 0 15916 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_165
timestamp 1
transform 1 0 16284 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_169
timestamp 1
transform 1 0 16652 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_177
timestamp 1
transform 1 0 17388 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_184
timestamp 1
transform 1 0 18032 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_202
timestamp 1
transform 1 0 19688 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_212
timestamp 1562078211
transform 1 0 20608 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_225
timestamp 1562078211
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_237
timestamp 1562078211
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_249
timestamp 1562078211
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_261
timestamp 1562078211
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_273
timestamp 1
transform 1 0 26220 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_277
timestamp 1
transform 1 0 26588 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_281
timestamp 1562078211
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_293
timestamp 1
transform 1 0 28060 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_297
timestamp 1
transform 1 0 28428 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_3
timestamp 1562078211
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_15
timestamp 1562078211
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_76_29
timestamp 1
transform 1 0 3772 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_33
timestamp 1
transform 1 0 4140 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_35
timestamp 1
transform 1 0 4324 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_52
timestamp 1562078211
transform 1 0 5888 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_64
timestamp 1
transform 1 0 6992 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_81
timestamp 1
transform 1 0 8556 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_85
timestamp 1
transform 1 0 8924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_87
timestamp 1
transform 1 0 9108 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_93
timestamp 1
transform 1 0 9660 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_111
timestamp 1
transform 1 0 11316 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_121
timestamp 1
transform 1 0 12236 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_76_129
timestamp 1
transform 1 0 12972 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_141
timestamp 1
transform 1 0 14076 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_149
timestamp 1
transform 1 0 14812 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_167
timestamp 1
transform 1 0 16468 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_177
timestamp 1
transform 1 0 17388 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_183
timestamp 1
transform 1 0 17940 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_193
timestamp 1
transform 1 0 18860 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_197
timestamp 1
transform 1 0 19228 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_204
timestamp 1
transform 1 0 19872 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_211
timestamp 1
transform 1 0 20516 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_216
timestamp 1
transform 1 0 20976 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_220
timestamp 1562078211
transform 1 0 21344 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_232
timestamp 1562078211
transform 1 0 22448 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_76_244
timestamp 1
transform 1 0 23552 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_253
timestamp 1562078211
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_265
timestamp 1562078211
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_277
timestamp 1562078211
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_76_289
timestamp 1
transform 1 0 27692 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_297
timestamp 1
transform 1 0 28428 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_3
timestamp 1562078211
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_15
timestamp 1562078211
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_77_27
timestamp 1
transform 1 0 3588 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_35
timestamp 1
transform 1 0 4324 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_42
timestamp 1562078211
transform 1 0 4968 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_64
timestamp 1
transform 1 0 6992 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_77_82
timestamp 1
transform 1 0 8648 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_93
timestamp 1
transform 1 0 9660 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_113
timestamp 1
transform 1 0 11500 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_121
timestamp 1
transform 1 0 12236 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_123
timestamp 1
transform 1 0 12420 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_130
timestamp 1
transform 1 0 13064 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_139
timestamp 1
transform 1 0 13892 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_144
timestamp 1
transform 1 0 14352 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_146
timestamp 1
transform 1 0 14536 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_77_156
timestamp 1
transform 1 0 15456 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_160
timestamp 1
transform 1 0 15824 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_169
timestamp 1
transform 1 0 16652 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_178
timestamp 1
transform 1 0 17480 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_180
timestamp 1
transform 1 0 17664 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_197
timestamp 1
transform 1 0 19228 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_207
timestamp 1
transform 1 0 20148 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_213
timestamp 1
transform 1 0 20700 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_77_217
timestamp 1
transform 1 0 21068 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_221
timestamp 1
transform 1 0 21436 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_225
timestamp 1562078211
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_237
timestamp 1562078211
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_249
timestamp 1562078211
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_261
timestamp 1562078211
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_77_273
timestamp 1
transform 1 0 26220 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_277
timestamp 1
transform 1 0 26588 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_281
timestamp 1562078211
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_77_293
timestamp 1
transform 1 0 28060 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_297
timestamp 1
transform 1 0 28428 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_3
timestamp 1562078211
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_15
timestamp 1562078211
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_29
timestamp 1562078211
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_41
timestamp 1562078211
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_78_53
timestamp 1
transform 1 0 5980 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_61
timestamp 1
transform 1 0 6716 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_71
timestamp 1
transform 1 0 7636 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_78
timestamp 1
transform 1 0 8280 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_82
timestamp 1
transform 1 0 8648 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_78_85
timestamp 1
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_93
timestamp 1
transform 1 0 9660 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_100
timestamp 1
transform 1 0 10304 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_111
timestamp 1
transform 1 0 11316 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_121
timestamp 1
transform 1 0 12236 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_78_131
timestamp 1
transform 1 0 13156 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_141
timestamp 1
transform 1 0 14076 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_158
timestamp 1
transform 1 0 15640 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_78_168
timestamp 1
transform 1 0 16560 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_172
timestamp 1
transform 1 0 16928 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_78_190
timestamp 1
transform 1 0 18584 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_194
timestamp 1
transform 1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_197
timestamp 1
transform 1 0 19228 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_206
timestamp 1562078211
transform 1 0 20056 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_218
timestamp 1562078211
transform 1 0 21160 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_230
timestamp 1562078211
transform 1 0 22264 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_78_242
timestamp 1
transform 1 0 23368 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_253
timestamp 1562078211
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_265
timestamp 1562078211
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_277
timestamp 1562078211
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_78_289
timestamp 1
transform 1 0 27692 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_297
timestamp 1
transform 1 0 28428 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_3
timestamp 1562078211
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_15
timestamp 1562078211
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_27
timestamp 1562078211
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_39
timestamp 1562078211
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_79_51
timestamp 1
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_57
timestamp 1562078211
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_69
timestamp 1562078211
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_81
timestamp 1562078211
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_79_93
timestamp 1
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_101
timestamp 1
transform 1 0 10396 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_79_108
timestamp 1
transform 1 0 11040 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_113
timestamp 1
transform 1 0 11500 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_119
timestamp 1562078211
transform 1 0 12052 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_79_131
timestamp 1
transform 1 0 13156 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_135
timestamp 1
transform 1 0 13524 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_79_141
timestamp 1
transform 1 0 14076 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_148
timestamp 1
transform 1 0 14720 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_79_152
timestamp 1
transform 1 0 15088 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_163
timestamp 1
transform 1 0 16100 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_79_169
timestamp 1
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_179
timestamp 1
transform 1 0 17572 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_79_189
timestamp 1
transform 1 0 18492 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_197
timestamp 1
transform 1 0 19228 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_79_215
timestamp 1
transform 1 0 20884 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_225
timestamp 1562078211
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_237
timestamp 1562078211
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_249
timestamp 1562078211
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_261
timestamp 1562078211
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_79_273
timestamp 1
transform 1 0 26220 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_277
timestamp 1
transform 1 0 26588 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_281
timestamp 1562078211
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_79_293
timestamp 1
transform 1 0 28060 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_297
timestamp 1
transform 1 0 28428 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_3
timestamp 1562078211
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_15
timestamp 1562078211
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_29
timestamp 1562078211
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_41
timestamp 1562078211
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_53
timestamp 1562078211
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_65
timestamp 1562078211
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_77
timestamp 1
transform 1 0 8188 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_81
timestamp 1
transform 1 0 8556 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_85
timestamp 1562078211
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_97
timestamp 1562078211
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_109
timestamp 1562078211
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_121
timestamp 1562078211
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_133
timestamp 1
transform 1 0 13340 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_137
timestamp 1
transform 1 0 13708 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_141
timestamp 1562078211
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_153
timestamp 1562078211
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_165
timestamp 1562078211
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_177
timestamp 1562078211
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_189
timestamp 1
transform 1 0 18492 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_193
timestamp 1
transform 1 0 18860 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_197
timestamp 1562078211
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_209
timestamp 1562078211
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_221
timestamp 1562078211
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_233
timestamp 1562078211
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_245
timestamp 1
transform 1 0 23644 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_249
timestamp 1
transform 1 0 24012 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_253
timestamp 1562078211
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_265
timestamp 1562078211
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_277
timestamp 1562078211
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_80_289
timestamp 1
transform 1 0 27692 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_297
timestamp 1
transform 1 0 28428 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_3
timestamp 1562078211
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_15
timestamp 1562078211
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_27
timestamp 1562078211
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_39
timestamp 1562078211
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_51
timestamp 1
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_57
timestamp 1562078211
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_69
timestamp 1562078211
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_81
timestamp 1562078211
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_93
timestamp 1562078211
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_105
timestamp 1
transform 1 0 10764 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_109
timestamp 1
transform 1 0 11132 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_113
timestamp 1562078211
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_125
timestamp 1562078211
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_137
timestamp 1562078211
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_149
timestamp 1562078211
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_161
timestamp 1
transform 1 0 15916 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_165
timestamp 1
transform 1 0 16284 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_169
timestamp 1562078211
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_181
timestamp 1562078211
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_193
timestamp 1562078211
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_205
timestamp 1562078211
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_217
timestamp 1
transform 1 0 21068 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_221
timestamp 1
transform 1 0 21436 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_225
timestamp 1562078211
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_237
timestamp 1562078211
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_249
timestamp 1562078211
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_261
timestamp 1562078211
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_273
timestamp 1
transform 1 0 26220 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_277
timestamp 1
transform 1 0 26588 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_281
timestamp 1562078211
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_293
timestamp 1
transform 1 0 28060 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_297
timestamp 1
transform 1 0 28428 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_3
timestamp 1562078211
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_15
timestamp 1562078211
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_29
timestamp 1562078211
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_82_41
timestamp 1
transform 1 0 4876 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_48
timestamp 1
transform 1 0 5520 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_82_52
timestamp 1
transform 1 0 5888 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_57
timestamp 1562078211
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_69
timestamp 1562078211
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_81
timestamp 1
transform 1 0 8556 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_85
timestamp 1562078211
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_97
timestamp 1562078211
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_109
timestamp 1
transform 1 0 11132 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_113
timestamp 1562078211
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_125
timestamp 1562078211
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_137
timestamp 1
transform 1 0 13708 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_141
timestamp 1562078211
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_153
timestamp 1562078211
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_165
timestamp 1
transform 1 0 16284 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_169
timestamp 1562078211
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_181
timestamp 1562078211
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_193
timestamp 1
transform 1 0 18860 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_197
timestamp 1562078211
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_209
timestamp 1562078211
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_221
timestamp 1
transform 1 0 21436 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_223
timestamp 1
transform 1 0 21620 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_225
timestamp 1
transform 1 0 21804 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_82_243
timestamp 1
transform 1 0 23460 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_258
timestamp 1562078211
transform 1 0 24840 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_82_270
timestamp 1
transform 1 0 25944 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_281
timestamp 1562078211
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_82_293
timestamp 1
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_297
timestamp 1
transform 1 0 28428 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform 1 0 11500 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 12696 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 12328 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 10120 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform 1 0 10304 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform 1 0 11500 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform 1 0 8096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 7728 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform 1 0 11592 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 11224 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform 1 0 10212 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 9568 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 7360 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform 1 0 6440 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform 1 0 7176 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform 1 0 6716 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 12328 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 6900 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 7084 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform 1 0 7268 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 8372 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 8280 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 10212 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 10856 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 6164 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 9752 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 7636 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform 1 0 6440 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform 1 0 8924 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform 1 0 6992 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 7636 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 6808 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform 1 0 9752 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform 1 0 7176 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 14996 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform 1 0 6440 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform -1 0 10120 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform 1 0 9016 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform -1 0 9292 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform -1 0 7636 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform -1 0 7176 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform -1 0 10212 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform 1 0 8004 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 11408 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform -1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform -1 0 11316 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform -1 0 10396 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform -1 0 6164 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform -1 0 7176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform 1 0 9844 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform 1 0 4968 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform 1 0 6256 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform -1 0 7176 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform 1 0 14168 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1
transform 1 0 15548 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1
transform -1 0 4508 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1
transform 1 0 7728 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1
transform -1 0 17112 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1
transform 1 0 24288 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1
transform -1 0 21436 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1
transform -1 0 20516 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1
transform 1 0 18216 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1
transform -1 0 20056 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1
transform -1 0 24012 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1
transform 1 0 22356 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1
transform -1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1
transform 1 0 25392 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1
transform 1 0 19412 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1
transform -1 0 18860 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1
transform 1 0 19320 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1
transform -1 0 19320 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1
transform 1 0 21804 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1
transform 1 0 24472 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1
transform -1 0 24196 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1
transform -1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1
transform -1 0 22172 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1
transform 1 0 20516 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1
transform -1 0 17480 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1
transform -1 0 17480 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1
transform 1 0 14996 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1
transform 1 0 22816 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1
transform -1 0 22632 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1
transform 1 0 20884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1
transform 1 0 15272 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1
transform -1 0 17480 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1
transform -1 0 18400 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1
transform -1 0 19596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1
transform 1 0 19320 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1
transform 1 0 19504 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1
transform 1 0 20700 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1
transform 1 0 19872 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1
transform -1 0 20056 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1
transform -1 0 17480 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1
transform -1 0 26496 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1
transform -1 0 25208 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1
transform -1 0 25208 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1
transform -1 0 18952 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1
transform 1 0 24472 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1
transform -1 0 24748 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1
transform -1 0 23920 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1
transform -1 0 18492 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1
transform 1 0 19320 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1
transform -1 0 19504 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1
transform -1 0 18952 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1
transform -1 0 16744 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1
transform 1 0 11500 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1
transform -1 0 13156 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1
transform -1 0 17480 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1
transform 1 0 19320 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1
transform 1 0 11592 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1
transform -1 0 12972 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1
transform -1 0 12328 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1
transform -1 0 14076 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1
transform 1 0 12420 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1
transform 1 0 8740 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1
transform -1 0 13432 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1
transform -1 0 14168 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1
transform 1 0 16744 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1
transform -1 0 16100 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1
transform 1 0 10212 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1
transform 1 0 10580 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1
transform 1 0 12788 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1
transform 1 0 15180 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1
transform -1 0 10764 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1
transform -1 0 15180 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1
transform -1 0 12696 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1
transform -1 0 14076 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1
transform 1 0 11592 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1
transform 1 0 20976 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1
transform 1 0 19596 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1
transform 1 0 24472 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1
transform -1 0 25208 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1
transform 1 0 15824 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1
transform -1 0 22908 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1
transform 1 0 24472 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1
transform 1 0 14444 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1
transform -1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1
transform 1 0 13156 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1
transform 1 0 23092 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1
transform -1 0 22356 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1
transform -1 0 21988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1
transform -1 0 20884 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1
transform 1 0 16744 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1
transform -1 0 16652 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1
transform -1 0 22816 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1
transform 1 0 20240 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1
transform 1 0 17848 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1
transform -1 0 17480 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1
transform 1 0 17664 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1
transform -1 0 17020 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1
transform 1 0 19136 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1
transform -1 0 19596 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 5244 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 1748 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 1748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1748 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 1748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1
transform -1 0 28520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output8
timestamp 1
transform 1 0 21988 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output9
timestamp 1
transform 1 0 27048 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output10
timestamp 1
transform 1 0 27048 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output11
timestamp 1
transform 1 0 27048 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_83
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_84
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_85
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_86
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_87
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_88
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_89
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_90
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_91
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_92
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_93
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_94
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_95
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_96
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_97
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_98
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_99
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_100
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_101
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_102
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_103
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_104
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_105
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_106
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_107
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_108
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_109
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_110
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_111
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_112
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_113
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_114
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_115
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_116
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_117
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_118
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_119
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_120
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_121
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_122
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_123
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_124
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_125
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_126
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_127
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_128
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_129
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_130
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_131
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_132
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_133
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_134
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_135
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_136
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_137
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1
transform -1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_138
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1
transform -1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_139
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1
transform -1 0 28888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_140
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1
transform -1 0 28888 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_141
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1
transform -1 0 28888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_142
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1
transform -1 0 28888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_143
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1
transform -1 0 28888 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_144
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1
transform -1 0 28888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_145
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1
transform -1 0 28888 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_146
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1
transform -1 0 28888 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_147
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1
transform -1 0 28888 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_148
timestamp 1
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1
transform -1 0 28888 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_149
timestamp 1
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1
transform -1 0 28888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_150
timestamp 1
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1
transform -1 0 28888 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_151
timestamp 1
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1
transform -1 0 28888 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_152
timestamp 1
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 1
transform -1 0 28888 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_153
timestamp 1
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 1
transform -1 0 28888 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_154
timestamp 1
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 1
transform -1 0 28888 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_155
timestamp 1
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 1
transform -1 0 28888 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_156
timestamp 1
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 1
transform -1 0 28888 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_157
timestamp 1
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 1
transform -1 0 28888 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_158
timestamp 1
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 1
transform -1 0 28888 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_159
timestamp 1
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 1
transform -1 0 28888 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_160
timestamp 1
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 1
transform -1 0 28888 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_161
timestamp 1
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 1
transform -1 0 28888 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_162
timestamp 1
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 1
transform -1 0 28888 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_163
timestamp 1
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 1
transform -1 0 28888 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_164
timestamp 1
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 1
transform -1 0 28888 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_165
timestamp 1
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 1
transform -1 0 28888 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_19
timestamp 1
transform 1 0 28244 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_20
timestamp 1
transform -1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_21
timestamp 1
transform -1 0 24840 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_22
timestamp 1
transform -1 0 1748 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_23
timestamp 1
transform -1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_24
timestamp 1
transform -1 0 1748 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_25
timestamp 1
transform -1 0 1748 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_26
timestamp 1
transform 1 0 28244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_27
timestamp 1
transform -1 0 1748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_28
timestamp 1
transform -1 0 28520 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_166
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_167
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_168
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_169
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_170
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_171
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_172
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_173
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_174
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_175
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_176
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_177
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_178
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_179
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_180
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_181
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_182
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_183
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_184
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_185
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_186
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_187
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_188
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_189
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_190
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_191
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_192
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_193
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_194
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_195
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_196
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_197
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_198
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_199
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_200
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_201
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_202
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_203
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_204
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_205
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_206
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_207
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_208
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_209
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_210
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_211
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_212
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_213
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_214
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_215
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_216
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_217
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_218
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_219
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_220
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_221
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_222
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_223
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_224
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_225
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_226
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_227
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_228
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_229
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_230
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_231
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_232
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_233
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_234
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_235
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_236
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_237
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_238
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_239
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_240
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_241
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_242
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_243
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_244
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_245
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_246
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_247
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_248
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_249
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_250
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_251
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_252
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_253
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_254
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_255
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_256
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_257
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_258
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_259
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_260
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_261
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_262
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_263
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_264
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_265
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_266
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_267
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_268
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_269
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_270
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_271
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_272
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_273
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_274
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_275
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_276
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_277
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_278
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_279
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_280
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_281
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_282
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_283
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_284
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_285
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_286
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_287
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_288
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_289
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_290
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_291
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_292
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_293
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_294
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_295
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_296
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_297
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_298
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_299
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_300
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_301
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_302
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_303
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_304
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_305
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_306
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_307
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_308
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_309
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_310
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_311
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_312
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_313
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_314
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_315
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_316
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_317
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_318
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_319
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_320
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_321
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_322
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_323
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_324
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_325
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_326
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_327
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_328
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_329
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_330
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_331
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_332
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_333
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_334
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_335
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_336
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_337
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_338
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_339
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_340
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_341
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_342
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_343
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_344
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_345
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_346
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_347
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_348
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_349
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_350
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_351
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_352
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_353
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_354
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_355
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_356
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_357
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_358
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_359
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_360
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_361
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_362
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_363
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_364
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_365
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_366
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_367
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_368
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_369
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_370
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_371
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_372
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_373
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_374
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_375
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_376
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_377
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_378
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_379
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_380
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_381
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_382
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_383
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_384
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_385
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_386
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_387
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_388
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_389
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_390
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_391
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_392
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_393
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_394
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_395
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_396
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_397
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_398
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_399
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_400
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_401
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_402
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_403
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_404
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_405
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_406
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_407
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_408
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_409
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_410
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_411
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_412
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_413
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_414
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_415
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_416
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_417
timestamp 1
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_418
timestamp 1
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_419
timestamp 1
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_420
timestamp 1
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_421
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_422
timestamp 1
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_423
timestamp 1
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_424
timestamp 1
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_425
timestamp 1
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_426
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_427
timestamp 1
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_428
timestamp 1
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_429
timestamp 1
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_430
timestamp 1
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_431
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_432
timestamp 1
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_433
timestamp 1
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_434
timestamp 1
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_435
timestamp 1
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_436
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_437
timestamp 1
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_438
timestamp 1
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_439
timestamp 1
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_440
timestamp 1
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_441
timestamp 1
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_442
timestamp 1
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_443
timestamp 1
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_444
timestamp 1
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_445
timestamp 1
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_446
timestamp 1
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_447
timestamp 1
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_448
timestamp 1
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_449
timestamp 1
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_450
timestamp 1
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_451
timestamp 1
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_452
timestamp 1
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_453
timestamp 1
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_454
timestamp 1
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_455
timestamp 1
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_456
timestamp 1
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_457
timestamp 1
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_458
timestamp 1
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_459
timestamp 1
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_460
timestamp 1
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_461
timestamp 1
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_462
timestamp 1
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_463
timestamp 1
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_464
timestamp 1
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_465
timestamp 1
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_466
timestamp 1
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_467
timestamp 1
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_468
timestamp 1
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_469
timestamp 1
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_470
timestamp 1
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_471
timestamp 1
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_472
timestamp 1
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_473
timestamp 1
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_474
timestamp 1
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_475
timestamp 1
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_476
timestamp 1
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_477
timestamp 1
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_478
timestamp 1
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_479
timestamp 1
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_480
timestamp 1
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_481
timestamp 1
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_482
timestamp 1
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_483
timestamp 1
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_484
timestamp 1
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_485
timestamp 1
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_486
timestamp 1
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_487
timestamp 1
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_488
timestamp 1
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_489
timestamp 1
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_490
timestamp 1
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_491
timestamp 1
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_492
timestamp 1
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_493
timestamp 1
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_494
timestamp 1
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_495
timestamp 1
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_496
timestamp 1
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_497
timestamp 1
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_498
timestamp 1
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_499
timestamp 1
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_500
timestamp 1
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_501
timestamp 1
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_502
timestamp 1
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_503
timestamp 1
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_504
timestamp 1
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_505
timestamp 1
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_506
timestamp 1
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_507
timestamp 1
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_508
timestamp 1
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_509
timestamp 1
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_510
timestamp 1
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_511
timestamp 1
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_512
timestamp 1
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_513
timestamp 1
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_514
timestamp 1
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_515
timestamp 1
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_516
timestamp 1
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_517
timestamp 1
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_518
timestamp 1
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_519
timestamp 1
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_520
timestamp 1
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_521
timestamp 1
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_522
timestamp 1
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_523
timestamp 1
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_524
timestamp 1
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_525
timestamp 1
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_526
timestamp 1
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_527
timestamp 1
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_528
timestamp 1
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_529
timestamp 1
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_530
timestamp 1
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_531
timestamp 1
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_532
timestamp 1
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_533
timestamp 1
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_534
timestamp 1
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_535
timestamp 1
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_536
timestamp 1
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_537
timestamp 1
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_538
timestamp 1
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_539
timestamp 1
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_540
timestamp 1
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_541
timestamp 1
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_542
timestamp 1
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_543
timestamp 1
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_544
timestamp 1
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_545
timestamp 1
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_546
timestamp 1
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_547
timestamp 1
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_548
timestamp 1
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_549
timestamp 1
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_550
timestamp 1
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_551
timestamp 1
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_552
timestamp 1
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_553
timestamp 1
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_554
timestamp 1
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_555
timestamp 1
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_556
timestamp 1
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_557
timestamp 1
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_558
timestamp 1
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_559
timestamp 1
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_560
timestamp 1
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_561
timestamp 1
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_562
timestamp 1
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_563
timestamp 1
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_564
timestamp 1
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_565
timestamp 1
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_566
timestamp 1
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_567
timestamp 1
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_568
timestamp 1
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_569
timestamp 1
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_570
timestamp 1
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_571
timestamp 1
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_572
timestamp 1
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_573
timestamp 1
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_574
timestamp 1
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_575
timestamp 1
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_576
timestamp 1
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_577
timestamp 1
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_578
timestamp 1
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_579
timestamp 1
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_580
timestamp 1
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_581
timestamp 1
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_582
timestamp 1
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_583
timestamp 1
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_584
timestamp 1
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_585
timestamp 1
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_586
timestamp 1
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_587
timestamp 1
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_588
timestamp 1
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_589
timestamp 1
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_590
timestamp 1
transform 1 0 26864 0 1 46784
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 5170 49200 5226 50000 0 FreeSans 224 90 0 0 enc0_a
port 1 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 enc0_b
port 2 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 enc1_a
port 3 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 enc1_b
port 4 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 enc2_a
port 5 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 enc2_b
port 6 nsew signal input
flabel metal3 s 29200 31288 30000 31408 0 FreeSans 480 0 0 0 io_oeb_high[0]
port 7 nsew signal output
flabel metal3 s 29200 27208 30000 27328 0 FreeSans 480 0 0 0 io_oeb_high[1]
port 8 nsew signal output
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 io_oeb_high[2]
port 9 nsew signal output
flabel metal2 s 24490 49200 24546 50000 0 FreeSans 224 90 0 0 io_oeb_high[3]
port 10 nsew signal output
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 io_oeb_high[4]
port 11 nsew signal output
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 io_oeb_high[5]
port 12 nsew signal output
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 io_oeb_low[0]
port 13 nsew signal output
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 io_oeb_low[1]
port 14 nsew signal output
flabel metal3 s 29200 14288 30000 14408 0 FreeSans 480 0 0 0 io_oeb_low[2]
port 15 nsew signal output
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 io_oeb_low[3]
port 16 nsew signal output
flabel metal2 s 21914 49200 21970 50000 0 FreeSans 224 90 0 0 pwm0_out
port 17 nsew signal output
flabel metal3 s 29200 31968 30000 32088 0 FreeSans 480 0 0 0 pwm1_out
port 18 nsew signal output
flabel metal3 s 29200 15648 30000 15768 0 FreeSans 480 0 0 0 pwm2_out
port 19 nsew signal output
flabel metal3 s 29200 8168 30000 8288 0 FreeSans 480 0 0 0 reset
port 20 nsew signal input
flabel metal3 s 29200 17008 30000 17128 0 FreeSans 480 0 0 0 sync
port 21 nsew signal output
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 22 nsew power bidirectional
flabel metal4 s 4868 2128 5188 47376 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 50000
<< end >>
