magic
tech sky130A
magscale 1 2
timestamp 1757431050
<< viali >>
rect 6745 47141 6779 47175
rect 6561 47005 6595 47039
rect 7113 45441 7147 45475
rect 11989 45441 12023 45475
rect 12265 45441 12299 45475
rect 6929 45373 6963 45407
rect 12081 45373 12115 45407
rect 7297 45237 7331 45271
rect 12173 45237 12207 45271
rect 12449 45237 12483 45271
rect 11621 45033 11655 45067
rect 13921 44965 13955 44999
rect 10241 44897 10275 44931
rect 12541 44897 12575 44931
rect 14197 44897 14231 44931
rect 14841 44897 14875 44931
rect 15301 44897 15335 44931
rect 7389 44829 7423 44863
rect 9505 44829 9539 44863
rect 12265 44829 12299 44863
rect 15117 44829 15151 44863
rect 7634 44761 7668 44795
rect 10508 44761 10542 44795
rect 12786 44761 12820 44795
rect 14933 44761 14967 44795
rect 8769 44693 8803 44727
rect 8953 44693 8987 44727
rect 11713 44693 11747 44727
rect 11253 44489 11287 44523
rect 12725 44489 12759 44523
rect 12817 44489 12851 44523
rect 13185 44489 13219 44523
rect 9045 44421 9079 44455
rect 10118 44421 10152 44455
rect 8309 44353 8343 44387
rect 8401 44353 8435 44387
rect 8861 44353 8895 44387
rect 9873 44353 9907 44387
rect 12357 44353 12391 44387
rect 12909 44353 12943 44387
rect 14309 44353 14343 44387
rect 14565 44353 14599 44387
rect 8677 44285 8711 44319
rect 9137 44285 9171 44319
rect 9781 44285 9815 44319
rect 12541 44285 12575 44319
rect 8585 44149 8619 44183
rect 11805 44149 11839 44183
rect 13093 44149 13127 44183
rect 11529 43945 11563 43979
rect 13093 43945 13127 43979
rect 13185 43945 13219 43979
rect 13277 43945 13311 43979
rect 10609 43877 10643 43911
rect 9229 43809 9263 43843
rect 11897 43809 11931 43843
rect 12265 43809 12299 43843
rect 12541 43809 12575 43843
rect 13553 43809 13587 43843
rect 9485 43741 9519 43775
rect 11713 43741 11747 43775
rect 12173 43741 12207 43775
rect 12633 43741 12667 43775
rect 13001 43741 13035 43775
rect 13461 43741 13495 43775
rect 13737 43741 13771 43775
rect 13921 43741 13955 43775
rect 14105 43741 14139 43775
rect 14657 43741 14691 43775
rect 11989 43673 12023 43707
rect 12449 43605 12483 43639
rect 12725 43605 12759 43639
rect 14105 43401 14139 43435
rect 11710 43265 11744 43299
rect 11805 43265 11839 43299
rect 12725 43265 12759 43299
rect 12992 43265 13026 43299
rect 19901 43265 19935 43299
rect 20168 43265 20202 43299
rect 12081 43197 12115 43231
rect 11529 43061 11563 43095
rect 12633 43061 12667 43095
rect 21281 43061 21315 43095
rect 12449 42857 12483 42891
rect 13093 42857 13127 42891
rect 11069 42721 11103 42755
rect 21649 42721 21683 42755
rect 11336 42653 11370 42687
rect 12541 42653 12575 42687
rect 12817 42653 12851 42687
rect 13277 42653 13311 42687
rect 13369 42653 13403 42687
rect 12633 42517 12667 42551
rect 13001 42517 13035 42551
rect 21097 42517 21131 42551
rect 13093 42177 13127 42211
rect 12541 41973 12575 42007
rect 20177 41769 20211 41803
rect 20269 41701 20303 41735
rect 20637 41701 20671 41735
rect 17141 41565 17175 41599
rect 20177 41565 20211 41599
rect 20637 41565 20671 41599
rect 20821 41565 20855 41599
rect 22845 41565 22879 41599
rect 26617 41565 26651 41599
rect 26801 41565 26835 41599
rect 16874 41497 16908 41531
rect 20545 41497 20579 41531
rect 23112 41497 23146 41531
rect 15761 41429 15795 41463
rect 20453 41429 20487 41463
rect 24225 41429 24259 41463
rect 26709 41429 26743 41463
rect 16681 41225 16715 41259
rect 23489 41225 23523 41259
rect 23765 41225 23799 41259
rect 17233 41157 17267 41191
rect 27230 41157 27264 41191
rect 16865 41089 16899 41123
rect 17417 41089 17451 41123
rect 17509 41089 17543 41123
rect 23397 41089 23431 41123
rect 23581 41089 23615 41123
rect 24133 41089 24167 41123
rect 26433 41089 26467 41123
rect 17141 41021 17175 41055
rect 24225 41021 24259 41055
rect 24409 41021 24443 41055
rect 26341 41021 26375 41055
rect 26985 41021 27019 41055
rect 17233 40953 17267 40987
rect 17049 40885 17083 40919
rect 26709 40885 26743 40919
rect 28365 40885 28399 40919
rect 20453 40681 20487 40715
rect 21097 40681 21131 40715
rect 23213 40681 23247 40715
rect 26709 40681 26743 40715
rect 20821 40545 20855 40579
rect 22937 40545 22971 40579
rect 23765 40545 23799 40579
rect 27169 40545 27203 40579
rect 27353 40545 27387 40579
rect 20637 40477 20671 40511
rect 20913 40477 20947 40511
rect 21005 40477 21039 40511
rect 21189 40477 21223 40511
rect 22845 40477 22879 40511
rect 23673 40477 23707 40511
rect 24409 40477 24443 40511
rect 26157 40477 26191 40511
rect 26341 40477 26375 40511
rect 26433 40477 26467 40511
rect 26617 40477 26651 40511
rect 27721 40477 27755 40511
rect 27997 40477 28031 40511
rect 23305 40341 23339 40375
rect 24501 40341 24535 40375
rect 26065 40341 26099 40375
rect 27077 40341 27111 40375
rect 27537 40341 27571 40375
rect 27905 40341 27939 40375
rect 21103 40137 21137 40171
rect 23397 40137 23431 40171
rect 23765 40137 23799 40171
rect 26985 40137 27019 40171
rect 27905 40137 27939 40171
rect 10609 40069 10643 40103
rect 21189 40069 21223 40103
rect 27445 40069 27479 40103
rect 27721 40069 27755 40103
rect 12081 40001 12115 40035
rect 12348 40001 12382 40035
rect 19809 40001 19843 40035
rect 19993 40001 20027 40035
rect 20637 40001 20671 40035
rect 20821 40001 20855 40035
rect 21005 40001 21039 40035
rect 21281 40001 21315 40035
rect 23213 40001 23247 40035
rect 23305 40001 23339 40035
rect 23949 40001 23983 40035
rect 24133 40001 24167 40035
rect 24409 40001 24443 40035
rect 24685 40001 24719 40035
rect 27537 40001 27571 40035
rect 9321 39933 9355 39967
rect 20913 39933 20947 39967
rect 23673 39933 23707 39967
rect 24041 39933 24075 39967
rect 24225 39933 24259 39967
rect 24869 39933 24903 39967
rect 27169 39865 27203 39899
rect 8769 39797 8803 39831
rect 13461 39797 13495 39831
rect 19993 39797 20027 39831
rect 20453 39797 20487 39831
rect 24501 39797 24535 39831
rect 10977 39593 11011 39627
rect 17601 39593 17635 39627
rect 18061 39593 18095 39627
rect 20269 39593 20303 39627
rect 21097 39593 21131 39627
rect 24133 39593 24167 39627
rect 12541 39457 12575 39491
rect 16773 39457 16807 39491
rect 20453 39457 20487 39491
rect 20729 39457 20763 39491
rect 21281 39457 21315 39491
rect 24777 39457 24811 39491
rect 8493 39389 8527 39423
rect 8585 39389 8619 39423
rect 8953 39389 8987 39423
rect 16865 39389 16899 39423
rect 17877 39389 17911 39423
rect 18245 39389 18279 39423
rect 19625 39389 19659 39423
rect 19809 39389 19843 39423
rect 19901 39389 19935 39423
rect 20085 39389 20119 39423
rect 20545 39389 20579 39423
rect 20637 39389 20671 39423
rect 21373 39389 21407 39423
rect 21649 39389 21683 39423
rect 23765 39389 23799 39423
rect 24041 39389 24075 39423
rect 24225 39389 24259 39423
rect 24593 39389 24627 39423
rect 8769 39321 8803 39355
rect 9198 39321 9232 39355
rect 12265 39321 12299 39355
rect 12808 39321 12842 39355
rect 17693 39321 17727 39355
rect 21741 39321 21775 39355
rect 23581 39321 23615 39355
rect 23949 39321 23983 39355
rect 10333 39253 10367 39287
rect 13921 39253 13955 39287
rect 17233 39253 17267 39287
rect 18337 39253 18371 39287
rect 19441 39253 19475 39287
rect 20913 39253 20947 39287
rect 24409 39253 24443 39287
rect 9045 39049 9079 39083
rect 13185 39049 13219 39083
rect 16221 39049 16255 39083
rect 18889 39049 18923 39083
rect 21005 39049 21039 39083
rect 19340 38981 19374 39015
rect 7665 38913 7699 38947
rect 7932 38913 7966 38947
rect 9597 38913 9631 38947
rect 9864 38913 9898 38947
rect 13369 38913 13403 38947
rect 13461 38913 13495 38947
rect 14565 38913 14599 38947
rect 14749 38913 14783 38947
rect 16037 38913 16071 38947
rect 16221 38913 16255 38947
rect 16313 38913 16347 38947
rect 16497 38913 16531 38947
rect 16681 38913 16715 38947
rect 16937 38913 16971 38947
rect 18337 38913 18371 38947
rect 18613 38913 18647 38947
rect 20913 38913 20947 38947
rect 23213 38913 23247 38947
rect 16405 38845 16439 38879
rect 18521 38845 18555 38879
rect 18889 38845 18923 38879
rect 19073 38845 19107 38879
rect 21189 38845 21223 38879
rect 23121 38845 23155 38879
rect 18061 38777 18095 38811
rect 20453 38777 20487 38811
rect 23581 38777 23615 38811
rect 10977 38709 11011 38743
rect 14657 38709 14691 38743
rect 18153 38709 18187 38743
rect 18705 38709 18739 38743
rect 20545 38709 20579 38743
rect 8125 38505 8159 38539
rect 9873 38505 9907 38539
rect 14289 38505 14323 38539
rect 15669 38505 15703 38539
rect 16773 38505 16807 38539
rect 16865 38505 16899 38539
rect 19533 38505 19567 38539
rect 20085 38505 20119 38539
rect 13921 38437 13955 38471
rect 14841 38437 14875 38471
rect 9505 38369 9539 38403
rect 10701 38369 10735 38403
rect 13461 38369 13495 38403
rect 17325 38369 17359 38403
rect 17417 38369 17451 38403
rect 19901 38369 19935 38403
rect 27169 38369 27203 38403
rect 8309 38301 8343 38335
rect 8493 38301 8527 38335
rect 9689 38301 9723 38335
rect 10609 38301 10643 38335
rect 11253 38301 11287 38335
rect 13553 38301 13587 38335
rect 14197 38301 14231 38335
rect 14565 38301 14599 38335
rect 14657 38301 14691 38335
rect 15393 38301 15427 38335
rect 15669 38301 15703 38335
rect 16589 38301 16623 38335
rect 16773 38301 16807 38335
rect 17693 38301 17727 38335
rect 17969 38301 18003 38335
rect 18245 38301 18279 38335
rect 19349 38301 19383 38335
rect 19533 38301 19567 38335
rect 19809 38301 19843 38335
rect 20545 38301 20579 38335
rect 27077 38301 27111 38335
rect 14933 38233 14967 38267
rect 15117 38233 15151 38267
rect 17785 38233 17819 38267
rect 18153 38233 18187 38267
rect 9965 38165 9999 38199
rect 15301 38165 15335 38199
rect 15485 38165 15519 38199
rect 17233 38165 17267 38199
rect 18337 38165 18371 38199
rect 20453 38165 20487 38199
rect 26709 38165 26743 38199
rect 8585 37961 8619 37995
rect 9781 37961 9815 37995
rect 17125 37961 17159 37995
rect 23765 37961 23799 37995
rect 26985 37961 27019 37995
rect 9505 37893 9539 37927
rect 9873 37893 9907 37927
rect 12449 37893 12483 37927
rect 17325 37893 17359 37927
rect 9229 37825 9263 37859
rect 9689 37825 9723 37859
rect 12265 37825 12299 37859
rect 12817 37825 12851 37859
rect 14105 37825 14139 37859
rect 14197 37825 14231 37859
rect 14289 37825 14323 37859
rect 14381 37825 14415 37859
rect 23673 37825 23707 37859
rect 27353 37825 27387 37859
rect 11161 37757 11195 37791
rect 12541 37757 12575 37791
rect 14565 37757 14599 37791
rect 23949 37757 23983 37791
rect 27261 37757 27295 37791
rect 10057 37621 10091 37655
rect 10609 37621 10643 37655
rect 16957 37621 16991 37655
rect 17141 37621 17175 37655
rect 23305 37621 23339 37655
rect 8953 37417 8987 37451
rect 10149 37417 10183 37451
rect 24501 37417 24535 37451
rect 8677 37349 8711 37383
rect 26801 37349 26835 37383
rect 27169 37349 27203 37383
rect 10333 37281 10367 37315
rect 7297 37213 7331 37247
rect 8953 37213 8987 37247
rect 9137 37213 9171 37247
rect 9229 37213 9263 37247
rect 10425 37213 10459 37247
rect 10701 37213 10735 37247
rect 12173 37213 12207 37247
rect 22845 37213 22879 37247
rect 24409 37213 24443 37247
rect 26709 37213 26743 37247
rect 26893 37213 26927 37247
rect 27077 37213 27111 37247
rect 27169 37213 27203 37247
rect 27353 37213 27387 37247
rect 27905 37213 27939 37247
rect 28457 37213 28491 37247
rect 7564 37145 7598 37179
rect 10149 37145 10183 37179
rect 10968 37145 11002 37179
rect 12440 37145 12474 37179
rect 23112 37145 23146 37179
rect 26617 37145 26651 37179
rect 9413 37077 9447 37111
rect 10609 37077 10643 37111
rect 12081 37077 12115 37111
rect 13553 37077 13587 37111
rect 24225 37077 24259 37111
rect 8033 36873 8067 36907
rect 9781 36873 9815 36907
rect 10885 36873 10919 36907
rect 12265 36873 12299 36907
rect 23213 36873 23247 36907
rect 26709 36873 26743 36907
rect 10517 36805 10551 36839
rect 10609 36805 10643 36839
rect 27230 36805 27264 36839
rect 8217 36737 8251 36771
rect 9597 36737 9631 36771
rect 10057 36737 10091 36771
rect 10333 36737 10367 36771
rect 10701 36737 10735 36771
rect 12449 36737 12483 36771
rect 12541 36737 12575 36771
rect 20913 36737 20947 36771
rect 23121 36737 23155 36771
rect 23305 36737 23339 36771
rect 26801 36737 26835 36771
rect 26985 36737 27019 36771
rect 8401 36669 8435 36703
rect 8861 36669 8895 36703
rect 9413 36669 9447 36703
rect 9689 36669 9723 36703
rect 9965 36669 9999 36703
rect 10241 36669 10275 36703
rect 28365 36533 28399 36567
rect 9505 36193 9539 36227
rect 22201 36193 22235 36227
rect 20453 36057 20487 36091
rect 8953 35989 8987 36023
rect 9321 35785 9355 35819
rect 9229 35717 9263 35751
rect 19533 35717 19567 35751
rect 6561 35649 6595 35683
rect 6837 35649 6871 35683
rect 7093 35649 7127 35683
rect 8953 35649 8987 35683
rect 9045 35649 9079 35683
rect 10445 35649 10479 35683
rect 19441 35649 19475 35683
rect 19717 35649 19751 35683
rect 28273 35649 28307 35683
rect 6377 35581 6411 35615
rect 6745 35581 6779 35615
rect 10701 35581 10735 35615
rect 26985 35581 27019 35615
rect 8217 35513 8251 35547
rect 19717 35445 19751 35479
rect 27629 35445 27663 35479
rect 28457 35445 28491 35479
rect 6377 35241 6411 35275
rect 11805 35241 11839 35275
rect 11897 35241 11931 35275
rect 28273 35241 28307 35275
rect 7021 35105 7055 35139
rect 12265 35105 12299 35139
rect 19533 35105 19567 35139
rect 11161 35037 11195 35071
rect 12081 35037 12115 35071
rect 19441 35037 19475 35071
rect 19717 35037 19751 35071
rect 19809 35037 19843 35071
rect 19993 35037 20027 35071
rect 20085 35037 20119 35071
rect 20361 35037 20395 35071
rect 20913 35037 20947 35071
rect 26893 35037 26927 35071
rect 27160 35037 27194 35071
rect 8401 34969 8435 35003
rect 9321 34969 9355 35003
rect 20545 34969 20579 35003
rect 10609 34901 10643 34935
rect 20177 34901 20211 34935
rect 20729 34901 20763 34935
rect 6193 34697 6227 34731
rect 10701 34697 10735 34731
rect 20361 34697 20395 34731
rect 21649 34697 21683 34731
rect 24133 34697 24167 34731
rect 26433 34697 26467 34731
rect 9588 34629 9622 34663
rect 21373 34629 21407 34663
rect 23765 34629 23799 34663
rect 23857 34629 23891 34663
rect 24777 34629 24811 34663
rect 26801 34629 26835 34663
rect 27721 34629 27755 34663
rect 4813 34561 4847 34595
rect 5069 34561 5103 34595
rect 16230 34561 16264 34595
rect 18521 34561 18555 34595
rect 18613 34561 18647 34595
rect 18797 34561 18831 34595
rect 18889 34561 18923 34595
rect 21097 34561 21131 34595
rect 21281 34561 21315 34595
rect 21465 34561 21499 34595
rect 22017 34561 22051 34595
rect 22201 34561 22235 34595
rect 22293 34561 22327 34595
rect 22569 34561 22603 34595
rect 22753 34561 22787 34595
rect 23489 34561 23523 34595
rect 23582 34561 23616 34595
rect 23995 34561 24029 34595
rect 24593 34561 24627 34595
rect 26341 34561 26375 34595
rect 26709 34561 26743 34595
rect 26985 34561 27019 34595
rect 27169 34561 27203 34595
rect 27537 34561 27571 34595
rect 9321 34493 9355 34527
rect 16497 34493 16531 34527
rect 19625 34493 19659 34527
rect 20177 34493 20211 34527
rect 20913 34493 20947 34527
rect 22385 34493 22419 34527
rect 27261 34493 27295 34527
rect 27353 34493 27387 34527
rect 19073 34425 19107 34459
rect 26617 34425 26651 34459
rect 15117 34357 15151 34391
rect 24961 34357 24995 34391
rect 16221 34153 16255 34187
rect 23121 34153 23155 34187
rect 25789 34153 25823 34187
rect 18061 34085 18095 34119
rect 18429 34017 18463 34051
rect 18981 34017 19015 34051
rect 20637 34017 20671 34051
rect 21741 34017 21775 34051
rect 22845 34017 22879 34051
rect 27997 34017 28031 34051
rect 15761 33949 15795 33983
rect 16037 33949 16071 33983
rect 16221 33949 16255 33983
rect 17785 33949 17819 33983
rect 17969 33949 18003 33983
rect 18337 33949 18371 33983
rect 20729 33949 20763 33983
rect 21925 33949 21959 33983
rect 25237 33949 25271 33983
rect 25421 33949 25455 33983
rect 25605 33949 25639 33983
rect 15577 33881 15611 33915
rect 18061 33881 18095 33915
rect 18245 33881 18279 33915
rect 20370 33881 20404 33915
rect 22109 33881 22143 33915
rect 22937 33881 22971 33915
rect 25513 33881 25547 33915
rect 15945 33813 15979 33847
rect 17877 33813 17911 33847
rect 19257 33813 19291 33847
rect 22201 33813 22235 33847
rect 23137 33813 23171 33847
rect 23305 33813 23339 33847
rect 27445 33813 27479 33847
rect 3709 33609 3743 33643
rect 15945 33609 15979 33643
rect 16681 33609 16715 33643
rect 17049 33609 17083 33643
rect 17601 33609 17635 33643
rect 19165 33609 19199 33643
rect 21189 33609 21223 33643
rect 23213 33609 23247 33643
rect 15301 33541 15335 33575
rect 17141 33541 17175 33575
rect 18030 33541 18064 33575
rect 19441 33541 19475 33575
rect 19641 33541 19675 33575
rect 19901 33541 19935 33575
rect 3525 33473 3559 33507
rect 12808 33473 12842 33507
rect 15025 33473 15059 33507
rect 15120 33473 15154 33507
rect 15577 33473 15611 33507
rect 16497 33473 16531 33507
rect 17509 33473 17543 33507
rect 17785 33473 17819 33507
rect 22100 33473 22134 33507
rect 23305 33473 23339 33507
rect 23489 33473 23523 33507
rect 3341 33405 3375 33439
rect 12541 33405 12575 33439
rect 14565 33405 14599 33439
rect 15485 33405 15519 33439
rect 16037 33405 16071 33439
rect 17233 33405 17267 33439
rect 21833 33405 21867 33439
rect 13921 33337 13955 33371
rect 16129 33337 16163 33371
rect 14013 33269 14047 33303
rect 19625 33269 19659 33303
rect 19809 33269 19843 33303
rect 23305 33269 23339 33303
rect 1593 33065 1627 33099
rect 13277 33065 13311 33099
rect 13553 33065 13587 33099
rect 18521 33065 18555 33099
rect 21281 33065 21315 33099
rect 21649 33065 21683 33099
rect 23213 33065 23247 33099
rect 25237 33065 25271 33099
rect 25421 32997 25455 33031
rect 12357 32929 12391 32963
rect 12817 32929 12851 32963
rect 12909 32929 12943 32963
rect 18429 32929 18463 32963
rect 21005 32929 21039 32963
rect 21833 32929 21867 32963
rect 23857 32929 23891 32963
rect 24869 32929 24903 32963
rect 27629 32929 27663 32963
rect 28181 32929 28215 32963
rect 1409 32861 1443 32895
rect 12265 32861 12299 32895
rect 12449 32861 12483 32895
rect 12541 32861 12575 32895
rect 12725 32861 12759 32895
rect 13093 32861 13127 32895
rect 15301 32861 15335 32895
rect 15393 32861 15427 32895
rect 15577 32861 15611 32895
rect 18705 32861 18739 32895
rect 21189 32861 21223 32895
rect 21465 32861 21499 32895
rect 24041 32861 24075 32895
rect 24225 32861 24259 32895
rect 24685 32861 24719 32895
rect 26617 32861 26651 32895
rect 26709 32861 26743 32895
rect 26985 32861 27019 32895
rect 13737 32793 13771 32827
rect 20738 32793 20772 32827
rect 22100 32793 22134 32827
rect 24133 32793 24167 32827
rect 25053 32793 25087 32827
rect 26893 32793 26927 32827
rect 13369 32725 13403 32759
rect 13537 32725 13571 32759
rect 15761 32725 15795 32759
rect 18889 32725 18923 32759
rect 19625 32725 19659 32759
rect 23305 32725 23339 32759
rect 24501 32725 24535 32759
rect 25253 32725 25287 32759
rect 26794 32725 26828 32759
rect 27169 32725 27203 32759
rect 12633 32521 12667 32555
rect 13461 32521 13495 32555
rect 19901 32521 19935 32555
rect 20729 32521 20763 32555
rect 22201 32521 22235 32555
rect 25053 32521 25087 32555
rect 26525 32521 26559 32555
rect 28365 32521 28399 32555
rect 12173 32385 12207 32419
rect 13001 32385 13035 32419
rect 13553 32385 13587 32419
rect 13737 32385 13771 32419
rect 14013 32385 14047 32419
rect 14105 32385 14139 32419
rect 14197 32385 14231 32419
rect 14381 32385 14415 32419
rect 14657 32385 14691 32419
rect 19257 32385 19291 32419
rect 20729 32385 20763 32419
rect 20821 32385 20855 32419
rect 21005 32385 21039 32419
rect 22385 32385 22419 32419
rect 22569 32385 22603 32419
rect 22661 32385 22695 32419
rect 23673 32385 23707 32419
rect 23940 32385 23974 32419
rect 25145 32385 25179 32419
rect 25412 32385 25446 32419
rect 26985 32385 27019 32419
rect 27241 32385 27275 32419
rect 12265 32317 12299 32351
rect 13093 32317 13127 32351
rect 13185 32317 13219 32351
rect 13277 32317 13311 32351
rect 14565 32249 14599 32283
rect 1409 32181 1443 32215
rect 11989 32181 12023 32215
rect 13921 32181 13955 32215
rect 14749 32181 14783 32215
rect 13001 31977 13035 32011
rect 14105 31977 14139 32011
rect 24409 31977 24443 32011
rect 24777 31977 24811 32011
rect 26617 31977 26651 32011
rect 26985 31977 27019 32011
rect 11805 31909 11839 31943
rect 28457 31909 28491 31943
rect 12817 31841 12851 31875
rect 13369 31841 13403 31875
rect 24133 31841 24167 31875
rect 25513 31841 25547 31875
rect 26341 31841 26375 31875
rect 26525 31841 26559 31875
rect 1409 31773 1443 31807
rect 8953 31773 8987 31807
rect 11713 31773 11747 31807
rect 11897 31773 11931 31807
rect 12541 31773 12575 31807
rect 13277 31773 13311 31807
rect 13921 31773 13955 31807
rect 14289 31773 14323 31807
rect 14381 31773 14415 31807
rect 24041 31773 24075 31807
rect 24225 31773 24259 31807
rect 24593 31773 24627 31807
rect 24869 31773 24903 31807
rect 24961 31773 24995 31807
rect 26801 31773 26835 31807
rect 28273 31773 28307 31807
rect 9198 31705 9232 31739
rect 13553 31705 13587 31739
rect 13737 31705 13771 31739
rect 10333 31637 10367 31671
rect 25789 31637 25823 31671
rect 8677 31433 8711 31467
rect 13553 31433 13587 31467
rect 25421 31433 25455 31467
rect 13369 31365 13403 31399
rect 25605 31365 25639 31399
rect 5641 31297 5675 31331
rect 6561 31297 6595 31331
rect 8493 31297 8527 31331
rect 11805 31297 11839 31331
rect 11897 31297 11931 31331
rect 11989 31297 12023 31331
rect 12173 31297 12207 31331
rect 12817 31297 12851 31331
rect 13185 31297 13219 31331
rect 24961 31297 24995 31331
rect 25053 31297 25087 31331
rect 25237 31297 25271 31331
rect 25513 31297 25547 31331
rect 25697 31297 25731 31331
rect 5825 31229 5859 31263
rect 6745 31229 6779 31263
rect 8309 31229 8343 31263
rect 8769 31229 8803 31263
rect 9321 31229 9355 31263
rect 13093 31229 13127 31263
rect 5457 31093 5491 31127
rect 6377 31093 6411 31127
rect 11529 31093 11563 31127
rect 6469 30889 6503 30923
rect 12817 30889 12851 30923
rect 1409 30753 1443 30787
rect 5273 30753 5307 30787
rect 5733 30753 5767 30787
rect 7113 30753 7147 30787
rect 7205 30753 7239 30787
rect 15669 30753 15703 30787
rect 5457 30685 5491 30719
rect 6377 30685 6411 30719
rect 7481 30685 7515 30719
rect 11253 30685 11287 30719
rect 11520 30685 11554 30719
rect 12725 30685 12759 30719
rect 12909 30685 12943 30719
rect 15577 30685 15611 30719
rect 7573 30617 7607 30651
rect 5641 30549 5675 30583
rect 7389 30549 7423 30583
rect 7757 30549 7791 30583
rect 12633 30549 12667 30583
rect 15945 30549 15979 30583
rect 6644 30277 6678 30311
rect 15761 30277 15795 30311
rect 5080 30209 5114 30243
rect 6377 30209 6411 30243
rect 9985 30209 10019 30243
rect 10241 30209 10275 30243
rect 10517 30209 10551 30243
rect 15301 30209 15335 30243
rect 15853 30209 15887 30243
rect 16313 30209 16347 30243
rect 16497 30209 16531 30243
rect 26985 30209 27019 30243
rect 27241 30209 27275 30243
rect 4813 30141 4847 30175
rect 8401 30141 8435 30175
rect 10333 30141 10367 30175
rect 10701 30141 10735 30175
rect 15209 30141 15243 30175
rect 15669 30141 15703 30175
rect 16129 30141 16163 30175
rect 7757 30073 7791 30107
rect 16037 30073 16071 30107
rect 16313 30073 16347 30107
rect 28365 30073 28399 30107
rect 6193 30005 6227 30039
rect 7849 30005 7883 30039
rect 8861 30005 8895 30039
rect 16221 30005 16255 30039
rect 5273 29801 5307 29835
rect 6837 29801 6871 29835
rect 11345 29801 11379 29835
rect 1593 29733 1627 29767
rect 6745 29733 6779 29767
rect 8769 29733 8803 29767
rect 6929 29665 6963 29699
rect 7389 29665 7423 29699
rect 8953 29665 8987 29699
rect 9321 29665 9355 29699
rect 10241 29665 10275 29699
rect 17049 29665 17083 29699
rect 1409 29597 1443 29631
rect 2973 29597 3007 29631
rect 3065 29597 3099 29631
rect 3893 29597 3927 29631
rect 5365 29597 5399 29631
rect 7113 29597 7147 29631
rect 9413 29597 9447 29631
rect 10425 29597 10459 29631
rect 11253 29597 11287 29631
rect 16782 29597 16816 29631
rect 3249 29529 3283 29563
rect 4138 29529 4172 29563
rect 5632 29529 5666 29563
rect 6837 29529 6871 29563
rect 7645 29529 7679 29563
rect 9045 29529 9079 29563
rect 7297 29461 7331 29495
rect 9229 29461 9263 29495
rect 9597 29461 9631 29495
rect 9689 29461 9723 29495
rect 11069 29461 11103 29495
rect 15669 29461 15703 29495
rect 5549 29257 5583 29291
rect 7573 29257 7607 29291
rect 10241 29257 10275 29291
rect 8769 29189 8803 29223
rect 9106 29189 9140 29223
rect 6193 29121 6227 29155
rect 7297 29121 7331 29155
rect 7389 29121 7423 29155
rect 8493 29121 8527 29155
rect 8585 29121 8619 29155
rect 8861 29121 8895 29155
rect 10333 29121 10367 29155
rect 10517 29121 10551 29155
rect 10609 29121 10643 29155
rect 15117 29121 15151 29155
rect 18337 29121 18371 29155
rect 18429 29121 18463 29155
rect 18613 29121 18647 29155
rect 1409 28985 1443 29019
rect 15209 28985 15243 29019
rect 18613 28985 18647 29019
rect 10333 28917 10367 28951
rect 10793 28917 10827 28951
rect 18429 28713 18463 28747
rect 21189 28645 21223 28679
rect 18061 28577 18095 28611
rect 9137 28509 9171 28543
rect 9505 28509 9539 28543
rect 17785 28509 17819 28543
rect 17877 28509 17911 28543
rect 18153 28509 18187 28543
rect 18245 28509 18279 28543
rect 18338 28509 18372 28543
rect 19809 28509 19843 28543
rect 19993 28509 20027 28543
rect 20913 28509 20947 28543
rect 21189 28509 21223 28543
rect 9229 28441 9263 28475
rect 9321 28441 9355 28475
rect 8953 28373 8987 28407
rect 17601 28373 17635 28407
rect 19901 28373 19935 28407
rect 21005 28373 21039 28407
rect 18153 28169 18187 28203
rect 19441 28169 19475 28203
rect 17877 28101 17911 28135
rect 20576 28101 20610 28135
rect 17509 28033 17543 28067
rect 17602 28033 17636 28067
rect 17785 28033 17819 28067
rect 18015 28033 18049 28067
rect 20821 28033 20855 28067
rect 20913 27965 20947 27999
rect 28549 27897 28583 27931
rect 21557 27829 21591 27863
rect 16957 27557 16991 27591
rect 18153 27557 18187 27591
rect 21465 27557 21499 27591
rect 22201 27557 22235 27591
rect 21557 27489 21591 27523
rect 22017 27489 22051 27523
rect 22109 27489 22143 27523
rect 13461 27421 13495 27455
rect 13645 27421 13679 27455
rect 17601 27421 17635 27455
rect 17877 27421 17911 27455
rect 17969 27421 18003 27455
rect 18797 27421 18831 27455
rect 18981 27421 19015 27455
rect 19073 27421 19107 27455
rect 19349 27421 19383 27455
rect 20821 27421 20855 27455
rect 21649 27421 21683 27455
rect 21833 27421 21867 27455
rect 22385 27421 22419 27455
rect 16681 27353 16715 27387
rect 17785 27353 17819 27387
rect 18613 27353 18647 27387
rect 19594 27353 19628 27387
rect 22569 27353 22603 27387
rect 13645 27285 13679 27319
rect 17141 27285 17175 27319
rect 20729 27285 20763 27319
rect 13185 27081 13219 27115
rect 17693 27081 17727 27115
rect 19073 27081 19107 27115
rect 9198 27013 9232 27047
rect 17509 27013 17543 27047
rect 20944 27013 20978 27047
rect 12725 26945 12759 26979
rect 13553 26945 13587 26979
rect 13829 26945 13863 26979
rect 14013 26945 14047 26979
rect 14105 26945 14139 26979
rect 14197 26945 14231 26979
rect 17325 26945 17359 26979
rect 19625 26945 19659 26979
rect 21189 26945 21223 26979
rect 8953 26877 8987 26911
rect 12633 26877 12667 26911
rect 13369 26877 13403 26911
rect 13461 26877 13495 26911
rect 13645 26877 13679 26911
rect 19809 26809 19843 26843
rect 10333 26741 10367 26775
rect 13093 26741 13127 26775
rect 14473 26741 14507 26775
rect 13461 26537 13495 26571
rect 15761 26537 15795 26571
rect 16681 26537 16715 26571
rect 19993 26537 20027 26571
rect 20453 26537 20487 26571
rect 13369 26469 13403 26503
rect 13829 26469 13863 26503
rect 19717 26469 19751 26503
rect 11989 26401 12023 26435
rect 13645 26333 13679 26367
rect 13921 26333 13955 26367
rect 14381 26333 14415 26367
rect 14637 26333 14671 26367
rect 17969 26333 18003 26367
rect 19349 26333 19383 26367
rect 19533 26333 19567 26367
rect 20269 26333 20303 26367
rect 20453 26333 20487 26367
rect 12256 26265 12290 26299
rect 19809 26265 19843 26299
rect 20009 26265 20043 26299
rect 20177 26197 20211 26231
rect 9229 25993 9263 26027
rect 12265 25993 12299 26027
rect 13553 25993 13587 26027
rect 16681 25993 16715 26027
rect 13921 25925 13955 25959
rect 16957 25925 16991 25959
rect 17049 25925 17083 25959
rect 17969 25925 18003 25959
rect 9413 25857 9447 25891
rect 9597 25857 9631 25891
rect 11989 25857 12023 25891
rect 12541 25857 12575 25891
rect 12633 25857 12667 25891
rect 12725 25857 12759 25891
rect 12909 25857 12943 25891
rect 13185 25857 13219 25891
rect 13645 25857 13679 25891
rect 16129 25857 16163 25891
rect 16221 25857 16255 25891
rect 16313 25857 16347 25891
rect 16860 25857 16894 25891
rect 17232 25857 17266 25891
rect 17325 25857 17359 25891
rect 17877 25857 17911 25891
rect 18183 25857 18217 25891
rect 18337 25857 18371 25891
rect 11805 25789 11839 25823
rect 13093 25789 13127 25823
rect 13921 25789 13955 25823
rect 17417 25789 17451 25823
rect 17601 25721 17635 25755
rect 12173 25653 12207 25687
rect 13737 25653 13771 25687
rect 15945 25653 15979 25687
rect 12449 25449 12483 25483
rect 13001 25381 13035 25415
rect 13277 25381 13311 25415
rect 6837 25313 6871 25347
rect 7021 25245 7055 25279
rect 12265 25245 12299 25279
rect 12449 25245 12483 25279
rect 12541 25245 12575 25279
rect 12817 25245 12851 25279
rect 13093 25245 13127 25279
rect 16037 25245 16071 25279
rect 16221 25245 16255 25279
rect 6592 25177 6626 25211
rect 12633 25177 12667 25211
rect 5457 25109 5491 25143
rect 7573 25109 7607 25143
rect 16129 25109 16163 25143
rect 13737 24905 13771 24939
rect 9036 24837 9070 24871
rect 1409 24769 1443 24803
rect 2697 24769 2731 24803
rect 3157 24769 3191 24803
rect 3424 24769 3458 24803
rect 4721 24769 4755 24803
rect 4977 24769 5011 24803
rect 7490 24769 7524 24803
rect 13553 24769 13587 24803
rect 13921 24769 13955 24803
rect 2513 24701 2547 24735
rect 2881 24701 2915 24735
rect 7757 24701 7791 24735
rect 8769 24701 8803 24735
rect 1593 24633 1627 24667
rect 14013 24633 14047 24667
rect 4537 24565 4571 24599
rect 6101 24565 6135 24599
rect 6377 24565 6411 24599
rect 10149 24565 10183 24599
rect 4813 24361 4847 24395
rect 7297 24361 7331 24395
rect 7849 24361 7883 24395
rect 13277 24293 13311 24327
rect 4445 24225 4479 24259
rect 4905 24225 4939 24259
rect 5457 24225 5491 24259
rect 6561 24225 6595 24259
rect 7389 24225 7423 24259
rect 13553 24225 13587 24259
rect 4629 24157 4663 24191
rect 6377 24157 6411 24191
rect 7573 24157 7607 24191
rect 8033 24157 8067 24191
rect 8125 24157 8159 24191
rect 13645 24157 13679 24191
rect 7297 24089 7331 24123
rect 5825 24021 5859 24055
rect 7205 24021 7239 24055
rect 7757 24021 7791 24055
rect 6561 23817 6595 23851
rect 7481 23817 7515 23851
rect 16313 23817 16347 23851
rect 17233 23817 17267 23851
rect 19257 23817 19291 23851
rect 6469 23749 6503 23783
rect 10241 23749 10275 23783
rect 15945 23749 15979 23783
rect 16037 23749 16071 23783
rect 16865 23749 16899 23783
rect 19409 23749 19443 23783
rect 19625 23749 19659 23783
rect 5917 23681 5951 23715
rect 6009 23681 6043 23715
rect 6745 23681 6779 23715
rect 7205 23681 7239 23715
rect 7297 23681 7331 23715
rect 9781 23681 9815 23715
rect 10425 23681 10459 23715
rect 15025 23681 15059 23715
rect 15301 23681 15335 23715
rect 15393 23681 15427 23715
rect 15669 23681 15703 23715
rect 15762 23681 15796 23715
rect 16134 23681 16168 23715
rect 16681 23681 16715 23715
rect 16957 23681 16991 23715
rect 17049 23681 17083 23715
rect 19717 23681 19751 23715
rect 19901 23681 19935 23715
rect 28273 23681 28307 23715
rect 6377 23613 6411 23647
rect 6837 23613 6871 23647
rect 9873 23613 9907 23647
rect 15577 23613 15611 23647
rect 10149 23545 10183 23579
rect 5733 23477 5767 23511
rect 7021 23477 7055 23511
rect 10609 23477 10643 23511
rect 15117 23477 15151 23511
rect 19441 23477 19475 23511
rect 19717 23477 19751 23511
rect 28457 23477 28491 23511
rect 10333 23273 10367 23307
rect 11437 23273 11471 23307
rect 16865 23273 16899 23307
rect 27721 23273 27755 23307
rect 12081 23205 12115 23239
rect 17049 23205 17083 23239
rect 5273 23137 5307 23171
rect 10701 23137 10735 23171
rect 10793 23137 10827 23171
rect 17417 23137 17451 23171
rect 18981 23137 19015 23171
rect 19993 23137 20027 23171
rect 20545 23137 20579 23171
rect 6745 23069 6779 23103
rect 7113 23069 7147 23103
rect 7389 23069 7423 23103
rect 8953 23069 8987 23103
rect 10425 23069 10459 23103
rect 11161 23069 11195 23103
rect 11253 23069 11287 23103
rect 11437 23069 11471 23103
rect 12173 23069 12207 23103
rect 17141 23069 17175 23103
rect 17233 23069 17267 23103
rect 18705 23069 18739 23103
rect 18889 23069 18923 23103
rect 19809 23069 19843 23103
rect 27537 23069 27571 23103
rect 5540 23001 5574 23035
rect 6929 23001 6963 23035
rect 7021 23001 7055 23035
rect 7656 23001 7690 23035
rect 9198 23001 9232 23035
rect 10910 23001 10944 23035
rect 11713 23001 11747 23035
rect 11897 23001 11931 23035
rect 16681 23001 16715 23035
rect 6653 22933 6687 22967
rect 7297 22933 7331 22967
rect 8769 22933 8803 22967
rect 11069 22933 11103 22967
rect 12357 22933 12391 22967
rect 16881 22933 16915 22967
rect 17141 22933 17175 22967
rect 18521 22933 18555 22967
rect 19257 22933 19291 22967
rect 6377 22729 6411 22763
rect 6745 22729 6779 22763
rect 8125 22729 8159 22763
rect 10609 22729 10643 22763
rect 14749 22729 14783 22763
rect 16221 22729 16255 22763
rect 19717 22729 19751 22763
rect 6561 22661 6595 22695
rect 8677 22661 8711 22695
rect 6653 22593 6687 22627
rect 6929 22593 6963 22627
rect 7481 22593 7515 22627
rect 8861 22593 8895 22627
rect 8953 22593 8987 22627
rect 9873 22593 9907 22627
rect 9965 22593 9999 22627
rect 10057 22593 10091 22627
rect 10149 22593 10183 22627
rect 10425 22593 10459 22627
rect 10609 22593 10643 22627
rect 14657 22593 14691 22627
rect 16129 22593 16163 22627
rect 16405 22593 16439 22627
rect 16681 22593 16715 22627
rect 17233 22593 17267 22627
rect 17693 22593 17727 22627
rect 17969 22593 18003 22627
rect 18245 22593 18279 22627
rect 18512 22593 18546 22627
rect 20830 22593 20864 22627
rect 21097 22593 21131 22627
rect 10333 22525 10367 22559
rect 17785 22525 17819 22559
rect 28549 22525 28583 22559
rect 16405 22457 16439 22491
rect 19625 22457 19659 22491
rect 18153 22389 18187 22423
rect 7297 22185 7331 22219
rect 11805 22185 11839 22219
rect 12817 22185 12851 22219
rect 18705 22185 18739 22219
rect 7113 22117 7147 22151
rect 6929 22049 6963 22083
rect 11713 22049 11747 22083
rect 18337 22049 18371 22083
rect 7297 21981 7331 22015
rect 7389 21981 7423 22015
rect 7573 21981 7607 22015
rect 11989 21981 12023 22015
rect 12173 21981 12207 22015
rect 12449 21981 12483 22015
rect 12633 21981 12667 22015
rect 12725 21981 12759 22015
rect 12817 21981 12851 22015
rect 12909 21981 12943 22015
rect 17150 21981 17184 22015
rect 17417 21981 17451 22015
rect 18521 21981 18555 22015
rect 18797 21981 18831 22015
rect 18981 21981 19015 22015
rect 12265 21913 12299 21947
rect 18889 21913 18923 21947
rect 6377 21845 6411 21879
rect 13185 21845 13219 21879
rect 16037 21845 16071 21879
rect 12633 21573 12667 21607
rect 12357 21369 12391 21403
rect 12173 21301 12207 21335
rect 7573 21097 7607 21131
rect 7021 20893 7055 20927
rect 12817 20893 12851 20927
rect 13001 20893 13035 20927
rect 7849 20825 7883 20859
rect 13001 20757 13035 20791
rect 9505 20485 9539 20519
rect 5917 20417 5951 20451
rect 6101 20417 6135 20451
rect 12081 20417 12115 20451
rect 12817 20417 12851 20451
rect 12909 20417 12943 20451
rect 13001 20417 13035 20451
rect 13185 20417 13219 20451
rect 14482 20417 14516 20451
rect 14749 20417 14783 20451
rect 14841 20417 14875 20451
rect 14933 20417 14967 20451
rect 15117 20417 15151 20451
rect 15853 20417 15887 20451
rect 16037 20417 16071 20451
rect 16129 20417 16163 20451
rect 12173 20349 12207 20383
rect 12449 20281 12483 20315
rect 5733 20213 5767 20247
rect 8217 20213 8251 20247
rect 12541 20213 12575 20247
rect 13369 20213 13403 20247
rect 15117 20213 15151 20247
rect 15853 20213 15887 20247
rect 6837 20009 6871 20043
rect 14197 20009 14231 20043
rect 14565 20009 14599 20043
rect 16681 20009 16715 20043
rect 13829 19941 13863 19975
rect 5457 19873 5491 19907
rect 14105 19873 14139 19907
rect 15301 19873 15335 19907
rect 17325 19873 17359 19907
rect 7481 19805 7515 19839
rect 12449 19805 12483 19839
rect 12705 19805 12739 19839
rect 14381 19805 14415 19839
rect 28549 19805 28583 19839
rect 5724 19737 5758 19771
rect 15568 19737 15602 19771
rect 6929 19669 6963 19703
rect 16773 19669 16807 19703
rect 6193 19465 6227 19499
rect 6377 19465 6411 19499
rect 7389 19465 7423 19499
rect 15669 19465 15703 19499
rect 6837 19397 6871 19431
rect 4813 19329 4847 19363
rect 5080 19329 5114 19363
rect 6561 19329 6595 19363
rect 7021 19329 7055 19363
rect 7481 19329 7515 19363
rect 15853 19329 15887 19363
rect 16037 19329 16071 19363
rect 16129 19329 16163 19363
rect 6745 19261 6779 19295
rect 7205 19261 7239 19295
rect 9597 19261 9631 19295
rect 8953 19125 8987 19159
rect 6745 18921 6779 18955
rect 23397 18853 23431 18887
rect 5365 18785 5399 18819
rect 8953 18785 8987 18819
rect 21373 18785 21407 18819
rect 5632 18717 5666 18751
rect 19533 18717 19567 18751
rect 21005 18717 21039 18751
rect 21189 18717 21223 18751
rect 21465 18717 21499 18751
rect 21649 18717 21683 18751
rect 22937 18717 22971 18751
rect 23029 18717 23063 18751
rect 23581 18717 23615 18751
rect 23765 18717 23799 18751
rect 23949 18717 23983 18751
rect 9198 18649 9232 18683
rect 19778 18649 19812 18683
rect 21557 18649 21591 18683
rect 10333 18581 10367 18615
rect 20913 18581 20947 18615
rect 23213 18581 23247 18615
rect 23857 18581 23891 18615
rect 9045 18377 9079 18411
rect 23397 18377 23431 18411
rect 8769 18241 8803 18275
rect 8881 18241 8915 18275
rect 10250 18241 10284 18275
rect 15209 18241 15243 18275
rect 15393 18241 15427 18275
rect 15761 18241 15795 18275
rect 16313 18241 16347 18275
rect 17969 18241 18003 18275
rect 20177 18241 20211 18275
rect 20444 18241 20478 18275
rect 22017 18241 22051 18275
rect 22284 18241 22318 18275
rect 23489 18241 23523 18275
rect 23756 18241 23790 18275
rect 25228 18241 25262 18275
rect 10517 18173 10551 18207
rect 24961 18173 24995 18207
rect 9137 18037 9171 18071
rect 15209 18037 15243 18071
rect 19257 18037 19291 18071
rect 21557 18037 21591 18071
rect 24869 18037 24903 18071
rect 26341 18037 26375 18071
rect 16037 17833 16071 17867
rect 19625 17833 19659 17867
rect 22385 17833 22419 17867
rect 23857 17833 23891 17867
rect 24041 17833 24075 17867
rect 25145 17833 25179 17867
rect 19993 17765 20027 17799
rect 22753 17765 22787 17799
rect 25513 17765 25547 17799
rect 20269 17697 20303 17731
rect 21833 17697 21867 17731
rect 23673 17697 23707 17731
rect 25605 17697 25639 17731
rect 26709 17697 26743 17731
rect 10149 17629 10183 17663
rect 10333 17629 10367 17663
rect 14657 17629 14691 17663
rect 18705 17629 18739 17663
rect 18797 17629 18831 17663
rect 19809 17629 19843 17663
rect 20085 17629 20119 17663
rect 20177 17629 20211 17663
rect 20361 17629 20395 17663
rect 21097 17629 21131 17663
rect 22569 17629 22603 17663
rect 22845 17629 22879 17663
rect 23121 17629 23155 17663
rect 24961 17629 24995 17663
rect 25329 17629 25363 17663
rect 26525 17629 26559 17663
rect 27261 17629 27295 17663
rect 14924 17561 14958 17595
rect 18521 17561 18555 17595
rect 20545 17561 20579 17595
rect 24009 17561 24043 17595
rect 24225 17561 24259 17595
rect 9965 17493 9999 17527
rect 18797 17493 18831 17527
rect 21281 17493 21315 17527
rect 24409 17493 24443 17527
rect 25973 17493 26007 17527
rect 20545 17289 20579 17323
rect 21297 17289 21331 17323
rect 21465 17289 21499 17323
rect 23029 17289 23063 17323
rect 23673 17289 23707 17323
rect 25605 17289 25639 17323
rect 18604 17221 18638 17255
rect 21097 17221 21131 17255
rect 11089 17153 11123 17187
rect 11345 17153 11379 17187
rect 16957 17153 16991 17187
rect 17141 17153 17175 17187
rect 17601 17153 17635 17187
rect 18337 17153 18371 17187
rect 20729 17153 20763 17187
rect 20913 17153 20947 17187
rect 21005 17153 21039 17187
rect 22937 17153 22971 17187
rect 23121 17153 23155 17187
rect 23213 17153 23247 17187
rect 23489 17153 23523 17187
rect 25421 17153 25455 17187
rect 25697 17153 25731 17187
rect 18245 17085 18279 17119
rect 20361 17085 20395 17119
rect 23305 17085 23339 17119
rect 19717 17017 19751 17051
rect 25421 17017 25455 17051
rect 9965 16949 9999 16983
rect 16957 16949 16991 16983
rect 19809 16949 19843 16983
rect 21281 16949 21315 16983
rect 9321 16745 9355 16779
rect 11529 16745 11563 16779
rect 12173 16745 12207 16779
rect 18429 16745 18463 16779
rect 18705 16745 18739 16779
rect 25605 16745 25639 16779
rect 10793 16677 10827 16711
rect 18889 16677 18923 16711
rect 25513 16677 25547 16711
rect 9505 16609 9539 16643
rect 10149 16609 10183 16643
rect 16589 16609 16623 16643
rect 26157 16609 26191 16643
rect 26893 16609 26927 16643
rect 6285 16541 6319 16575
rect 7757 16541 7791 16575
rect 9597 16541 9631 16575
rect 9873 16541 9907 16575
rect 9965 16541 9999 16575
rect 10885 16541 10919 16575
rect 11253 16541 11287 16575
rect 11713 16541 11747 16575
rect 11805 16541 11839 16575
rect 12357 16541 12391 16575
rect 12541 16541 12575 16575
rect 16856 16541 16890 16575
rect 18153 16541 18187 16575
rect 18429 16541 18463 16575
rect 25513 16541 25547 16575
rect 25881 16541 25915 16575
rect 11069 16473 11103 16507
rect 11161 16473 11195 16507
rect 18521 16473 18555 16507
rect 26801 16473 26835 16507
rect 27138 16473 27172 16507
rect 5733 16405 5767 16439
rect 7113 16405 7147 16439
rect 9689 16405 9723 16439
rect 11437 16405 11471 16439
rect 17969 16405 18003 16439
rect 18245 16405 18279 16439
rect 18721 16405 18755 16439
rect 25789 16405 25823 16439
rect 28273 16405 28307 16439
rect 5549 16201 5583 16235
rect 6193 16201 6227 16235
rect 7757 16201 7791 16235
rect 10609 16201 10643 16235
rect 11345 16201 11379 16235
rect 18981 16201 19015 16235
rect 25237 16201 25271 16235
rect 28457 16201 28491 16235
rect 6622 16133 6656 16167
rect 8217 16133 8251 16167
rect 12326 16133 12360 16167
rect 19165 16133 19199 16167
rect 24041 16133 24075 16167
rect 1409 16065 1443 16099
rect 4169 16065 4203 16099
rect 4425 16065 4459 16099
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 6377 16065 6411 16099
rect 10241 16065 10275 16099
rect 10333 16065 10367 16099
rect 10425 16065 10459 16099
rect 17794 16065 17828 16099
rect 18061 16065 18095 16099
rect 18889 16065 18923 16099
rect 23305 16065 23339 16099
rect 23489 16065 23523 16099
rect 23673 16065 23707 16099
rect 23857 16065 23891 16099
rect 24409 16065 24443 16099
rect 24685 16065 24719 16099
rect 24961 16065 24995 16099
rect 25053 16065 25087 16099
rect 28273 16065 28307 16099
rect 10701 15997 10735 16031
rect 12081 15997 12115 16031
rect 18705 15997 18739 16031
rect 23581 15997 23615 16031
rect 24225 15997 24259 16031
rect 24593 15997 24627 16031
rect 10057 15929 10091 15963
rect 24777 15929 24811 15963
rect 1593 15861 1627 15895
rect 9505 15861 9539 15895
rect 13461 15861 13495 15895
rect 16681 15861 16715 15895
rect 18153 15861 18187 15895
rect 19165 15861 19199 15895
rect 28181 15861 28215 15895
rect 3433 15657 3467 15691
rect 8309 15657 8343 15691
rect 11069 15657 11103 15691
rect 12633 15657 12667 15691
rect 17693 15657 17727 15691
rect 18153 15657 18187 15691
rect 3065 15521 3099 15555
rect 6285 15521 6319 15555
rect 8493 15521 8527 15555
rect 3249 15453 3283 15487
rect 6469 15453 6503 15487
rect 6745 15453 6779 15487
rect 8585 15453 8619 15487
rect 10517 15453 10551 15487
rect 11253 15453 11287 15487
rect 11520 15453 11554 15487
rect 17141 15453 17175 15487
rect 17785 15453 17819 15487
rect 17969 15453 18003 15487
rect 18245 15453 18279 15487
rect 19901 15453 19935 15487
rect 19994 15453 20028 15487
rect 20366 15453 20400 15487
rect 21465 15453 21499 15487
rect 21558 15453 21592 15487
rect 6653 15385 6687 15419
rect 6990 15385 7024 15419
rect 8309 15385 8343 15419
rect 8953 15385 8987 15419
rect 20177 15385 20211 15419
rect 20269 15385 20303 15419
rect 8125 15317 8159 15351
rect 8769 15317 8803 15351
rect 20545 15317 20579 15351
rect 21833 15317 21867 15351
rect 8677 15113 8711 15147
rect 10425 15113 10459 15147
rect 10977 15113 11011 15147
rect 22477 15113 22511 15147
rect 10517 15045 10551 15079
rect 14105 15045 14139 15079
rect 14289 15045 14323 15079
rect 14565 15045 14599 15079
rect 17693 15045 17727 15079
rect 22109 15045 22143 15079
rect 22201 15045 22235 15079
rect 7297 14977 7331 15011
rect 7564 14977 7598 15011
rect 9312 14977 9346 15011
rect 10793 14977 10827 15011
rect 13461 14977 13495 15011
rect 13921 14977 13955 15011
rect 14381 14977 14415 15011
rect 14657 14977 14691 15011
rect 14749 14977 14783 15011
rect 14933 14977 14967 15011
rect 17509 14977 17543 15011
rect 21925 14977 21959 15011
rect 22293 14977 22327 15011
rect 9045 14909 9079 14943
rect 10609 14909 10643 14943
rect 13553 14909 13587 14943
rect 14841 14909 14875 14943
rect 13829 14841 13863 14875
rect 10517 14773 10551 14807
rect 14381 14773 14415 14807
rect 17877 14773 17911 14807
rect 7665 14569 7699 14603
rect 9689 14569 9723 14603
rect 14197 14569 14231 14603
rect 18889 14569 18923 14603
rect 19809 14569 19843 14603
rect 20637 14501 20671 14535
rect 20821 14501 20855 14535
rect 8953 14433 8987 14467
rect 9597 14433 9631 14467
rect 10057 14433 10091 14467
rect 19349 14433 19383 14467
rect 7849 14365 7883 14399
rect 8033 14365 8067 14399
rect 8125 14365 8159 14399
rect 8677 14365 8711 14399
rect 9873 14365 9907 14399
rect 13461 14365 13495 14399
rect 13553 14365 13587 14399
rect 14105 14365 14139 14399
rect 14381 14365 14415 14399
rect 14565 14365 14599 14399
rect 16957 14365 16991 14399
rect 17049 14365 17083 14399
rect 17233 14365 17267 14399
rect 17325 14365 17359 14399
rect 18337 14365 18371 14399
rect 18613 14365 18647 14399
rect 18705 14365 18739 14399
rect 19257 14365 19291 14399
rect 19533 14365 19567 14399
rect 19625 14365 19659 14399
rect 13645 14297 13679 14331
rect 13737 14297 13771 14331
rect 17509 14297 17543 14331
rect 18521 14297 18555 14331
rect 21097 14297 21131 14331
rect 13921 14229 13955 14263
rect 14749 14229 14783 14263
rect 25605 14025 25639 14059
rect 18705 13957 18739 13991
rect 25145 13889 25179 13923
rect 25329 13889 25363 13923
rect 25697 13889 25731 13923
rect 24961 13821 24995 13855
rect 17233 13685 17267 13719
rect 24869 13685 24903 13719
rect 25053 13685 25087 13719
rect 13737 13481 13771 13515
rect 16313 13481 16347 13515
rect 24501 13481 24535 13515
rect 26157 13481 26191 13515
rect 12357 13345 12391 13379
rect 15393 13345 15427 13379
rect 24777 13345 24811 13379
rect 26801 13345 26835 13379
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 15577 13277 15611 13311
rect 15853 13277 15887 13311
rect 17141 13277 17175 13311
rect 21557 13277 21591 13311
rect 21741 13277 21775 13311
rect 24501 13277 24535 13311
rect 24685 13277 24719 13311
rect 25033 13277 25067 13311
rect 12624 13209 12658 13243
rect 16281 13209 16315 13243
rect 16497 13209 16531 13243
rect 26249 13209 26283 13243
rect 15669 13141 15703 13175
rect 16037 13141 16071 13175
rect 16129 13141 16163 13175
rect 21649 13141 21683 13175
rect 23213 12937 23247 12971
rect 23397 12937 23431 12971
rect 25237 12937 25271 12971
rect 16681 12869 16715 12903
rect 22078 12869 22112 12903
rect 17049 12801 17083 12835
rect 21281 12801 21315 12835
rect 21833 12801 21867 12835
rect 23305 12801 23339 12835
rect 24777 12801 24811 12835
rect 25605 12801 25639 12835
rect 16957 12733 16991 12767
rect 21373 12733 21407 12767
rect 24685 12733 24719 12767
rect 25513 12733 25547 12767
rect 17049 12665 17083 12699
rect 21649 12665 21683 12699
rect 25145 12665 25179 12699
rect 12633 12393 12667 12427
rect 16313 12393 16347 12427
rect 22017 12393 22051 12427
rect 23213 12325 23247 12359
rect 21465 12257 21499 12291
rect 22661 12257 22695 12291
rect 23305 12257 23339 12291
rect 9781 12189 9815 12223
rect 9965 12189 9999 12223
rect 12817 12189 12851 12223
rect 13001 12189 13035 12223
rect 16221 12189 16255 12223
rect 21557 12189 21591 12223
rect 22845 12189 22879 12223
rect 23029 12189 23063 12223
rect 22477 12121 22511 12155
rect 9597 12053 9631 12087
rect 21925 12053 21959 12087
rect 22385 12053 22419 12087
rect 15669 11849 15703 11883
rect 9404 11781 9438 11815
rect 16221 11781 16255 11815
rect 16773 11781 16807 11815
rect 15301 11713 15335 11747
rect 15485 11713 15519 11747
rect 15761 11713 15795 11747
rect 18429 11713 18463 11747
rect 9137 11645 9171 11679
rect 12081 11645 12115 11679
rect 17049 11645 17083 11679
rect 18521 11645 18555 11679
rect 16037 11577 16071 11611
rect 18061 11577 18095 11611
rect 10517 11509 10551 11543
rect 11529 11509 11563 11543
rect 15301 11509 15335 11543
rect 11713 11305 11747 11339
rect 13461 11305 13495 11339
rect 16313 11305 16347 11339
rect 21557 11305 21591 11339
rect 10333 11237 10367 11271
rect 15393 11237 15427 11271
rect 11069 11169 11103 11203
rect 12081 11169 12115 11203
rect 15117 11169 15151 11203
rect 15945 11169 15979 11203
rect 16037 11169 16071 11203
rect 22477 11169 22511 11203
rect 22569 11169 22603 11203
rect 22753 11169 22787 11203
rect 8953 11101 8987 11135
rect 15025 11101 15059 11135
rect 15853 11101 15887 11135
rect 16497 11101 16531 11135
rect 16589 11101 16623 11135
rect 21741 11101 21775 11135
rect 22109 11101 22143 11135
rect 22293 11101 22327 11135
rect 22385 11101 22419 11135
rect 9220 11033 9254 11067
rect 12348 11033 12382 11067
rect 21833 11033 21867 11067
rect 21925 11033 21959 11067
rect 15485 10965 15519 10999
rect 9413 10761 9447 10795
rect 12909 10761 12943 10795
rect 13185 10761 13219 10795
rect 15853 10761 15887 10795
rect 19901 10761 19935 10795
rect 24961 10761 24995 10795
rect 11805 10693 11839 10727
rect 13093 10693 13127 10727
rect 24593 10693 24627 10727
rect 25421 10693 25455 10727
rect 9597 10625 9631 10659
rect 11161 10625 11195 10659
rect 11345 10625 11379 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 14740 10625 14774 10659
rect 17969 10625 18003 10659
rect 18889 10625 18923 10659
rect 24501 10625 24535 10659
rect 24777 10625 24811 10659
rect 25053 10625 25087 10659
rect 25237 10625 25271 10659
rect 8769 10557 8803 10591
rect 9321 10557 9355 10591
rect 9781 10557 9815 10591
rect 12265 10557 12299 10591
rect 14473 10557 14507 10591
rect 18061 10557 18095 10591
rect 18797 10557 18831 10591
rect 19441 10557 19475 10591
rect 19533 10557 19567 10591
rect 19625 10557 19659 10591
rect 19717 10557 19751 10591
rect 12081 10489 12115 10523
rect 19257 10489 19291 10523
rect 10977 10421 11011 10455
rect 18245 10421 18279 10455
rect 10149 10217 10183 10251
rect 10609 10217 10643 10251
rect 11345 10217 11379 10251
rect 15209 10217 15243 10251
rect 24225 10217 24259 10251
rect 25697 10217 25731 10251
rect 11437 10149 11471 10183
rect 25145 10149 25179 10183
rect 11069 10081 11103 10115
rect 11161 10081 11195 10115
rect 17509 10081 17543 10115
rect 18429 10081 18463 10115
rect 18521 10081 18555 10115
rect 18889 10081 18923 10115
rect 19349 10081 19383 10115
rect 24501 10081 24535 10115
rect 25053 10081 25087 10115
rect 25513 10081 25547 10115
rect 1409 10013 1443 10047
rect 10333 10013 10367 10047
rect 10425 10013 10459 10047
rect 10701 10013 10735 10047
rect 12817 10013 12851 10047
rect 15025 10013 15059 10047
rect 15209 10013 15243 10047
rect 17693 10013 17727 10047
rect 18337 10013 18371 10047
rect 18797 10013 18831 10047
rect 19441 10013 19475 10047
rect 23949 10013 23983 10047
rect 24041 10013 24075 10047
rect 24593 10013 24627 10047
rect 25881 10013 25915 10047
rect 25973 10013 26007 10047
rect 10609 9945 10643 9979
rect 10793 9945 10827 9979
rect 12550 9945 12584 9979
rect 17877 9945 17911 9979
rect 10885 9877 10919 9911
rect 17969 9877 18003 9911
rect 19809 9877 19843 9911
rect 24961 9877 24995 9911
rect 26065 9877 26099 9911
rect 10333 9673 10367 9707
rect 10517 9673 10551 9707
rect 11529 9673 11563 9707
rect 18429 9673 18463 9707
rect 19441 9673 19475 9707
rect 25053 9673 25087 9707
rect 10241 9605 10275 9639
rect 14565 9605 14599 9639
rect 15025 9605 15059 9639
rect 15209 9605 15243 9639
rect 18797 9605 18831 9639
rect 24041 9605 24075 9639
rect 24409 9605 24443 9639
rect 25421 9605 25455 9639
rect 25605 9605 25639 9639
rect 7205 9537 7239 9571
rect 7461 9537 7495 9571
rect 9689 9537 9723 9571
rect 10149 9537 10183 9571
rect 10793 9537 10827 9571
rect 12642 9537 12676 9571
rect 14657 9537 14691 9571
rect 15301 9537 15335 9571
rect 18337 9537 18371 9571
rect 18613 9537 18647 9571
rect 19073 9537 19107 9571
rect 19257 9537 19291 9571
rect 21281 9537 21315 9571
rect 22017 9537 22051 9571
rect 23765 9537 23799 9571
rect 23949 9537 23983 9571
rect 24961 9537 24995 9571
rect 9505 9469 9539 9503
rect 12909 9469 12943 9503
rect 18981 9469 19015 9503
rect 21189 9469 21223 9503
rect 21649 9469 21683 9503
rect 21925 9469 21959 9503
rect 25145 9469 25179 9503
rect 8585 9401 8619 9435
rect 9965 9401 9999 9435
rect 24593 9401 24627 9435
rect 9873 9333 9907 9367
rect 11345 9333 11379 9367
rect 15025 9333 15059 9367
rect 22293 9333 22327 9367
rect 23949 9333 23983 9367
rect 9413 9129 9447 9163
rect 10517 9129 10551 9163
rect 10977 9129 11011 9163
rect 12173 9129 12207 9163
rect 15577 9129 15611 9163
rect 21741 9129 21775 9163
rect 25789 9129 25823 9163
rect 7205 9061 7239 9095
rect 22201 9061 22235 9095
rect 5825 8993 5859 9027
rect 8033 8993 8067 9027
rect 10609 8993 10643 9027
rect 12541 8993 12575 9027
rect 19717 8993 19751 9027
rect 19901 8993 19935 9027
rect 21649 8993 21683 9027
rect 24409 8993 24443 9027
rect 9965 8925 9999 8959
rect 10517 8925 10551 8959
rect 10793 8925 10827 8959
rect 11069 8925 11103 8959
rect 11713 8925 11747 8959
rect 11805 8925 11839 8959
rect 11989 8925 12023 8959
rect 14197 8925 14231 8959
rect 17233 8925 17267 8959
rect 17417 8925 17451 8959
rect 19625 8925 19659 8959
rect 20085 8925 20119 8959
rect 21925 8925 21959 8959
rect 22477 8925 22511 8959
rect 24665 8925 24699 8959
rect 6070 8857 6104 8891
rect 12357 8857 12391 8891
rect 14464 8857 14498 8891
rect 20177 8857 20211 8891
rect 22201 8857 22235 8891
rect 7481 8789 7515 8823
rect 17325 8789 17359 8823
rect 19257 8789 19291 8823
rect 22109 8789 22143 8823
rect 22385 8789 22419 8823
rect 5641 8585 5675 8619
rect 7297 8585 7331 8619
rect 10701 8585 10735 8619
rect 14749 8585 14783 8619
rect 18337 8585 18371 8619
rect 23213 8585 23247 8619
rect 28365 8585 28399 8619
rect 9588 8517 9622 8551
rect 11897 8517 11931 8551
rect 22100 8517 22134 8551
rect 5365 8449 5399 8483
rect 5457 8449 5491 8483
rect 7481 8449 7515 8483
rect 7573 8449 7607 8483
rect 10977 8449 11011 8483
rect 11161 8449 11195 8483
rect 14933 8449 14967 8483
rect 15209 8449 15243 8483
rect 16957 8449 16991 8483
rect 17224 8449 17258 8483
rect 18705 8449 18739 8483
rect 18889 8449 18923 8483
rect 21833 8449 21867 8483
rect 28549 8449 28583 8483
rect 9321 8381 9355 8415
rect 11713 8381 11747 8415
rect 15117 8381 15151 8415
rect 18889 8313 18923 8347
rect 10793 8245 10827 8279
rect 8953 8041 8987 8075
rect 20637 8041 20671 8075
rect 19257 7905 19291 7939
rect 10333 7837 10367 7871
rect 19513 7837 19547 7871
rect 10088 7769 10122 7803
rect 5457 2601 5491 2635
rect 5273 2397 5307 2431
rect 27169 2397 27203 2431
<< metal1 >>
rect 1104 47354 28888 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 28888 47354
rect 1104 47280 28888 47302
rect 6733 47175 6791 47181
rect 6733 47141 6745 47175
rect 6779 47172 6791 47175
rect 7098 47172 7104 47184
rect 6779 47144 7104 47172
rect 6779 47141 6791 47144
rect 6733 47135 6791 47141
rect 7098 47132 7104 47144
rect 7156 47132 7162 47184
rect 6546 46996 6552 47048
rect 6604 46996 6610 47048
rect 1104 46810 28888 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 28888 46810
rect 1104 46736 28888 46758
rect 1104 46266 28888 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 28888 46266
rect 1104 46192 28888 46214
rect 1104 45722 28888 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 28888 45722
rect 1104 45648 28888 45670
rect 7098 45432 7104 45484
rect 7156 45432 7162 45484
rect 11977 45475 12035 45481
rect 11977 45441 11989 45475
rect 12023 45441 12035 45475
rect 11977 45435 12035 45441
rect 12253 45475 12311 45481
rect 12253 45441 12265 45475
rect 12299 45472 12311 45475
rect 12342 45472 12348 45484
rect 12299 45444 12348 45472
rect 12299 45441 12311 45444
rect 12253 45435 12311 45441
rect 6917 45407 6975 45413
rect 6917 45373 6929 45407
rect 6963 45404 6975 45407
rect 8202 45404 8208 45416
rect 6963 45376 8208 45404
rect 6963 45373 6975 45376
rect 6917 45367 6975 45373
rect 8202 45364 8208 45376
rect 8260 45364 8266 45416
rect 11992 45336 12020 45435
rect 12342 45432 12348 45444
rect 12400 45432 12406 45484
rect 12066 45364 12072 45416
rect 12124 45364 12130 45416
rect 12250 45336 12256 45348
rect 11992 45308 12256 45336
rect 12250 45296 12256 45308
rect 12308 45296 12314 45348
rect 7282 45228 7288 45280
rect 7340 45228 7346 45280
rect 12158 45228 12164 45280
rect 12216 45228 12222 45280
rect 12434 45228 12440 45280
rect 12492 45228 12498 45280
rect 1104 45178 28888 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 28888 45178
rect 1104 45104 28888 45126
rect 11609 45067 11667 45073
rect 11609 45033 11621 45067
rect 11655 45064 11667 45067
rect 12066 45064 12072 45076
rect 11655 45036 12072 45064
rect 11655 45033 11667 45036
rect 11609 45027 11667 45033
rect 12066 45024 12072 45036
rect 12124 45024 12130 45076
rect 13909 44999 13967 45005
rect 13909 44965 13921 44999
rect 13955 44965 13967 44999
rect 13909 44959 13967 44965
rect 9582 44928 9588 44940
rect 9416 44900 9588 44928
rect 7377 44863 7435 44869
rect 7377 44829 7389 44863
rect 7423 44860 7435 44863
rect 9416 44860 9444 44900
rect 9582 44888 9588 44900
rect 9640 44928 9646 44940
rect 10229 44931 10287 44937
rect 10229 44928 10241 44931
rect 9640 44900 10241 44928
rect 9640 44888 9646 44900
rect 10229 44897 10241 44900
rect 10275 44897 10287 44931
rect 12526 44928 12532 44940
rect 10229 44891 10287 44897
rect 11256 44900 12532 44928
rect 7423 44832 9444 44860
rect 9493 44863 9551 44869
rect 7423 44829 7435 44832
rect 7377 44823 7435 44829
rect 9493 44829 9505 44863
rect 9539 44829 9551 44863
rect 10244 44860 10272 44891
rect 11256 44860 11284 44900
rect 12526 44888 12532 44900
rect 12584 44888 12590 44940
rect 13538 44888 13544 44940
rect 13596 44928 13602 44940
rect 13924 44928 13952 44959
rect 14185 44931 14243 44937
rect 14185 44928 14197 44931
rect 13596 44900 14197 44928
rect 13596 44888 13602 44900
rect 14185 44897 14197 44900
rect 14231 44897 14243 44931
rect 14185 44891 14243 44897
rect 14829 44931 14887 44937
rect 14829 44897 14841 44931
rect 14875 44928 14887 44931
rect 15289 44931 15347 44937
rect 15289 44928 15301 44931
rect 14875 44900 15301 44928
rect 14875 44897 14887 44900
rect 14829 44891 14887 44897
rect 15289 44897 15301 44900
rect 15335 44897 15347 44931
rect 15289 44891 15347 44897
rect 10244 44832 11284 44860
rect 9493 44823 9551 44829
rect 7282 44752 7288 44804
rect 7340 44792 7346 44804
rect 7622 44795 7680 44801
rect 7622 44792 7634 44795
rect 7340 44764 7634 44792
rect 7340 44752 7346 44764
rect 7622 44761 7634 44764
rect 7668 44761 7680 44795
rect 9508 44792 9536 44823
rect 12250 44820 12256 44872
rect 12308 44820 12314 44872
rect 13814 44820 13820 44872
rect 13872 44860 13878 44872
rect 15105 44863 15163 44869
rect 15105 44860 15117 44863
rect 13872 44832 15117 44860
rect 13872 44820 13878 44832
rect 15105 44829 15117 44832
rect 15151 44829 15163 44863
rect 15105 44823 15163 44829
rect 7622 44755 7680 44761
rect 8772 44764 9536 44792
rect 8772 44733 8800 44764
rect 8757 44727 8815 44733
rect 8757 44693 8769 44727
rect 8803 44693 8815 44727
rect 8757 44687 8815 44693
rect 8938 44684 8944 44736
rect 8996 44684 9002 44736
rect 9508 44724 9536 44764
rect 10496 44795 10554 44801
rect 10496 44761 10508 44795
rect 10542 44792 10554 44795
rect 11514 44792 11520 44804
rect 10542 44764 11520 44792
rect 10542 44761 10554 44764
rect 10496 44755 10554 44761
rect 11514 44752 11520 44764
rect 11572 44752 11578 44804
rect 12158 44792 12164 44804
rect 11624 44764 12164 44792
rect 11624 44724 11652 44764
rect 12158 44752 12164 44764
rect 12216 44752 12222 44804
rect 12618 44752 12624 44804
rect 12676 44792 12682 44804
rect 12774 44795 12832 44801
rect 12774 44792 12786 44795
rect 12676 44764 12786 44792
rect 12676 44752 12682 44764
rect 12774 44761 12786 44764
rect 12820 44761 12832 44795
rect 12774 44755 12832 44761
rect 14458 44752 14464 44804
rect 14516 44792 14522 44804
rect 14921 44795 14979 44801
rect 14921 44792 14933 44795
rect 14516 44764 14933 44792
rect 14516 44752 14522 44764
rect 14921 44761 14933 44764
rect 14967 44761 14979 44795
rect 14921 44755 14979 44761
rect 9508 44696 11652 44724
rect 11701 44727 11759 44733
rect 11701 44693 11713 44727
rect 11747 44724 11759 44727
rect 11882 44724 11888 44736
rect 11747 44696 11888 44724
rect 11747 44693 11759 44696
rect 11701 44687 11759 44693
rect 11882 44684 11888 44696
rect 11940 44684 11946 44736
rect 1104 44634 28888 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 28888 44634
rect 1104 44560 28888 44582
rect 11241 44523 11299 44529
rect 11241 44489 11253 44523
rect 11287 44520 11299 44523
rect 12250 44520 12256 44532
rect 11287 44492 12256 44520
rect 11287 44489 11299 44492
rect 11241 44483 11299 44489
rect 12250 44480 12256 44492
rect 12308 44520 12314 44532
rect 12713 44523 12771 44529
rect 12713 44520 12725 44523
rect 12308 44492 12725 44520
rect 12308 44480 12314 44492
rect 12713 44489 12725 44492
rect 12759 44489 12771 44523
rect 12713 44483 12771 44489
rect 12805 44523 12863 44529
rect 12805 44489 12817 44523
rect 12851 44520 12863 44523
rect 13173 44523 13231 44529
rect 13173 44520 13185 44523
rect 12851 44492 13185 44520
rect 12851 44489 12863 44492
rect 12805 44483 12863 44489
rect 13173 44489 13185 44492
rect 13219 44520 13231 44523
rect 13262 44520 13268 44532
rect 13219 44492 13268 44520
rect 13219 44489 13231 44492
rect 13173 44483 13231 44489
rect 13262 44480 13268 44492
rect 13320 44480 13326 44532
rect 8938 44452 8944 44464
rect 8312 44424 8944 44452
rect 8312 44393 8340 44424
rect 8938 44412 8944 44424
rect 8996 44412 9002 44464
rect 9033 44455 9091 44461
rect 9033 44421 9045 44455
rect 9079 44452 9091 44455
rect 10106 44455 10164 44461
rect 10106 44452 10118 44455
rect 9079 44424 10118 44452
rect 9079 44421 9091 44424
rect 9033 44415 9091 44421
rect 10106 44421 10118 44424
rect 10152 44421 10164 44455
rect 10106 44415 10164 44421
rect 12526 44412 12532 44464
rect 12584 44452 12590 44464
rect 12584 44424 14596 44452
rect 12584 44412 12590 44424
rect 8297 44387 8355 44393
rect 8297 44353 8309 44387
rect 8343 44353 8355 44387
rect 8297 44347 8355 44353
rect 8389 44387 8447 44393
rect 8389 44353 8401 44387
rect 8435 44384 8447 44387
rect 8849 44387 8907 44393
rect 8849 44384 8861 44387
rect 8435 44356 8861 44384
rect 8435 44353 8447 44356
rect 8389 44347 8447 44353
rect 8849 44353 8861 44356
rect 8895 44384 8907 44387
rect 8895 44356 9536 44384
rect 8895 44353 8907 44356
rect 8849 44347 8907 44353
rect 8665 44319 8723 44325
rect 8665 44285 8677 44319
rect 8711 44316 8723 44319
rect 9125 44319 9183 44325
rect 9125 44316 9137 44319
rect 8711 44288 9137 44316
rect 8711 44285 8723 44288
rect 8665 44279 8723 44285
rect 9125 44285 9137 44288
rect 9171 44285 9183 44319
rect 9125 44279 9183 44285
rect 9508 44248 9536 44356
rect 9582 44344 9588 44396
rect 9640 44384 9646 44396
rect 9861 44387 9919 44393
rect 9861 44384 9873 44387
rect 9640 44356 9873 44384
rect 9640 44344 9646 44356
rect 9861 44353 9873 44356
rect 9907 44353 9919 44387
rect 11698 44384 11704 44396
rect 9861 44347 9919 44353
rect 9968 44356 11704 44384
rect 9766 44276 9772 44328
rect 9824 44276 9830 44328
rect 9968 44316 9996 44356
rect 11698 44344 11704 44356
rect 11756 44344 11762 44396
rect 12066 44344 12072 44396
rect 12124 44384 12130 44396
rect 12345 44387 12403 44393
rect 12345 44384 12357 44387
rect 12124 44356 12357 44384
rect 12124 44344 12130 44356
rect 12345 44353 12357 44356
rect 12391 44384 12403 44387
rect 12897 44387 12955 44393
rect 12391 44356 12572 44384
rect 12391 44353 12403 44356
rect 12345 44347 12403 44353
rect 12544 44325 12572 44356
rect 12897 44353 12909 44387
rect 12943 44384 12955 44387
rect 13170 44384 13176 44396
rect 12943 44356 13176 44384
rect 12943 44353 12955 44356
rect 12897 44347 12955 44353
rect 13170 44344 13176 44356
rect 13228 44384 13234 44396
rect 13538 44384 13544 44396
rect 13228 44356 13544 44384
rect 13228 44344 13234 44356
rect 13538 44344 13544 44356
rect 13596 44344 13602 44396
rect 14297 44387 14355 44393
rect 14297 44353 14309 44387
rect 14343 44384 14355 44387
rect 14458 44384 14464 44396
rect 14343 44356 14464 44384
rect 14343 44353 14355 44356
rect 14297 44347 14355 44353
rect 14458 44344 14464 44356
rect 14516 44344 14522 44396
rect 14568 44393 14596 44424
rect 14553 44387 14611 44393
rect 14553 44353 14565 44387
rect 14599 44353 14611 44387
rect 14553 44347 14611 44353
rect 9876 44288 9996 44316
rect 12529 44319 12587 44325
rect 9876 44248 9904 44288
rect 12529 44285 12541 44319
rect 12575 44285 12587 44319
rect 12529 44279 12587 44285
rect 9508 44220 9904 44248
rect 8570 44140 8576 44192
rect 8628 44140 8634 44192
rect 11790 44140 11796 44192
rect 11848 44140 11854 44192
rect 12710 44140 12716 44192
rect 12768 44180 12774 44192
rect 13081 44183 13139 44189
rect 13081 44180 13093 44183
rect 12768 44152 13093 44180
rect 12768 44140 12774 44152
rect 13081 44149 13093 44152
rect 13127 44149 13139 44183
rect 13081 44143 13139 44149
rect 1104 44090 28888 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 28888 44090
rect 1104 44016 28888 44038
rect 9582 43976 9588 43988
rect 9232 43948 9588 43976
rect 9232 43849 9260 43948
rect 9582 43936 9588 43948
rect 9640 43936 9646 43988
rect 9858 43936 9864 43988
rect 9916 43976 9922 43988
rect 9916 43948 10640 43976
rect 9916 43936 9922 43948
rect 10612 43917 10640 43948
rect 11514 43936 11520 43988
rect 11572 43936 11578 43988
rect 12434 43936 12440 43988
rect 12492 43976 12498 43988
rect 13081 43979 13139 43985
rect 13081 43976 13093 43979
rect 12492 43948 13093 43976
rect 12492 43936 12498 43948
rect 13081 43945 13093 43948
rect 13127 43945 13139 43979
rect 13081 43939 13139 43945
rect 13170 43936 13176 43988
rect 13228 43936 13234 43988
rect 13262 43936 13268 43988
rect 13320 43936 13326 43988
rect 10597 43911 10655 43917
rect 10597 43877 10609 43911
rect 10643 43908 10655 43911
rect 12986 43908 12992 43920
rect 10643 43880 12296 43908
rect 10643 43877 10655 43880
rect 10597 43871 10655 43877
rect 9217 43843 9275 43849
rect 9217 43809 9229 43843
rect 9263 43809 9275 43843
rect 9217 43803 9275 43809
rect 11882 43800 11888 43852
rect 11940 43800 11946 43852
rect 12268 43849 12296 43880
rect 12452 43880 12992 43908
rect 12253 43843 12311 43849
rect 12253 43809 12265 43843
rect 12299 43840 12311 43843
rect 12342 43840 12348 43852
rect 12299 43812 12348 43840
rect 12299 43809 12311 43812
rect 12253 43803 12311 43809
rect 12342 43800 12348 43812
rect 12400 43800 12406 43852
rect 8570 43732 8576 43784
rect 8628 43772 8634 43784
rect 9473 43775 9531 43781
rect 9473 43772 9485 43775
rect 8628 43744 9485 43772
rect 8628 43732 8634 43744
rect 9473 43741 9485 43744
rect 9519 43741 9531 43775
rect 9473 43735 9531 43741
rect 11698 43732 11704 43784
rect 11756 43732 11762 43784
rect 12161 43775 12219 43781
rect 12161 43741 12173 43775
rect 12207 43772 12219 43775
rect 12452 43772 12480 43880
rect 12986 43868 12992 43880
rect 13044 43868 13050 43920
rect 12529 43843 12587 43849
rect 12529 43809 12541 43843
rect 12575 43840 12587 43843
rect 12710 43840 12716 43852
rect 12575 43812 12716 43840
rect 12575 43809 12587 43812
rect 12529 43803 12587 43809
rect 12710 43800 12716 43812
rect 12768 43800 12774 43852
rect 13541 43843 13599 43849
rect 13541 43840 13553 43843
rect 12912 43812 13553 43840
rect 12207 43744 12480 43772
rect 12207 43741 12219 43744
rect 12161 43735 12219 43741
rect 12618 43732 12624 43784
rect 12676 43772 12682 43784
rect 12912 43772 12940 43812
rect 13541 43809 13553 43812
rect 13587 43809 13599 43843
rect 13541 43803 13599 43809
rect 12676 43744 12940 43772
rect 12676 43732 12682 43744
rect 12986 43732 12992 43784
rect 13044 43772 13050 43784
rect 13170 43772 13176 43784
rect 13044 43744 13176 43772
rect 13044 43732 13050 43744
rect 13170 43732 13176 43744
rect 13228 43732 13234 43784
rect 13449 43775 13507 43781
rect 13449 43741 13461 43775
rect 13495 43741 13507 43775
rect 13449 43735 13507 43741
rect 13725 43775 13783 43781
rect 13725 43741 13737 43775
rect 13771 43772 13783 43775
rect 13814 43772 13820 43784
rect 13771 43744 13820 43772
rect 13771 43741 13783 43744
rect 13725 43735 13783 43741
rect 11977 43707 12035 43713
rect 11977 43673 11989 43707
rect 12023 43704 12035 43707
rect 13464 43704 13492 43735
rect 13814 43732 13820 43744
rect 13872 43732 13878 43784
rect 13909 43775 13967 43781
rect 13909 43741 13921 43775
rect 13955 43772 13967 43775
rect 14093 43775 14151 43781
rect 14093 43772 14105 43775
rect 13955 43744 14105 43772
rect 13955 43741 13967 43744
rect 13909 43735 13967 43741
rect 14093 43741 14105 43744
rect 14139 43741 14151 43775
rect 14093 43735 14151 43741
rect 14642 43732 14648 43784
rect 14700 43732 14706 43784
rect 14660 43704 14688 43732
rect 12023 43676 12664 43704
rect 13464 43676 14688 43704
rect 12023 43673 12035 43676
rect 11977 43667 12035 43673
rect 12636 43648 12664 43676
rect 12158 43596 12164 43648
rect 12216 43636 12222 43648
rect 12437 43639 12495 43645
rect 12437 43636 12449 43639
rect 12216 43608 12449 43636
rect 12216 43596 12222 43608
rect 12437 43605 12449 43608
rect 12483 43605 12495 43639
rect 12437 43599 12495 43605
rect 12618 43596 12624 43648
rect 12676 43596 12682 43648
rect 12713 43639 12771 43645
rect 12713 43605 12725 43639
rect 12759 43636 12771 43639
rect 12802 43636 12808 43648
rect 12759 43608 12808 43636
rect 12759 43605 12771 43608
rect 12713 43599 12771 43605
rect 12802 43596 12808 43608
rect 12860 43596 12866 43648
rect 1104 43546 28888 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 28888 43546
rect 1104 43472 28888 43494
rect 11698 43392 11704 43444
rect 11756 43432 11762 43444
rect 13354 43432 13360 43444
rect 11756 43404 13360 43432
rect 11756 43392 11762 43404
rect 13354 43392 13360 43404
rect 13412 43432 13418 43444
rect 13814 43432 13820 43444
rect 13412 43404 13820 43432
rect 13412 43392 13418 43404
rect 13814 43392 13820 43404
rect 13872 43392 13878 43444
rect 14093 43435 14151 43441
rect 14093 43401 14105 43435
rect 14139 43432 14151 43435
rect 14642 43432 14648 43444
rect 14139 43404 14648 43432
rect 14139 43401 14151 43404
rect 14093 43395 14151 43401
rect 14642 43392 14648 43404
rect 14700 43392 14706 43444
rect 22830 43364 22836 43376
rect 19904 43336 22836 43364
rect 11698 43296 11704 43308
rect 11659 43268 11704 43296
rect 11698 43256 11704 43268
rect 11756 43256 11762 43308
rect 11790 43256 11796 43308
rect 11848 43256 11854 43308
rect 12526 43256 12532 43308
rect 12584 43296 12590 43308
rect 12986 43305 12992 43308
rect 12713 43299 12771 43305
rect 12713 43296 12725 43299
rect 12584 43268 12725 43296
rect 12584 43256 12590 43268
rect 12713 43265 12725 43268
rect 12759 43265 12771 43299
rect 12713 43259 12771 43265
rect 12980 43259 12992 43305
rect 12986 43256 12992 43259
rect 13044 43256 13050 43308
rect 19904 43305 19932 43336
rect 22830 43324 22836 43336
rect 22888 43324 22894 43376
rect 20162 43305 20168 43308
rect 19889 43299 19947 43305
rect 19889 43265 19901 43299
rect 19935 43265 19947 43299
rect 19889 43259 19947 43265
rect 20156 43259 20168 43305
rect 20162 43256 20168 43259
rect 20220 43256 20226 43308
rect 12069 43231 12127 43237
rect 12069 43197 12081 43231
rect 12115 43228 12127 43231
rect 12434 43228 12440 43240
rect 12115 43200 12440 43228
rect 12115 43197 12127 43200
rect 12069 43191 12127 43197
rect 12434 43188 12440 43200
rect 12492 43188 12498 43240
rect 11330 43052 11336 43104
rect 11388 43092 11394 43104
rect 11517 43095 11575 43101
rect 11517 43092 11529 43095
rect 11388 43064 11529 43092
rect 11388 43052 11394 43064
rect 11517 43061 11529 43064
rect 11563 43061 11575 43095
rect 11517 43055 11575 43061
rect 12621 43095 12679 43101
rect 12621 43061 12633 43095
rect 12667 43092 12679 43095
rect 12710 43092 12716 43104
rect 12667 43064 12716 43092
rect 12667 43061 12679 43064
rect 12621 43055 12679 43061
rect 12710 43052 12716 43064
rect 12768 43052 12774 43104
rect 21266 43052 21272 43104
rect 21324 43052 21330 43104
rect 1104 43002 28888 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 28888 43002
rect 1104 42928 28888 42950
rect 12434 42848 12440 42900
rect 12492 42848 12498 42900
rect 12986 42848 12992 42900
rect 13044 42888 13050 42900
rect 13081 42891 13139 42897
rect 13081 42888 13093 42891
rect 13044 42860 13093 42888
rect 13044 42848 13050 42860
rect 13081 42857 13093 42860
rect 13127 42857 13139 42891
rect 13081 42851 13139 42857
rect 9582 42712 9588 42764
rect 9640 42752 9646 42764
rect 11057 42755 11115 42761
rect 11057 42752 11069 42755
rect 9640 42724 11069 42752
rect 9640 42712 9646 42724
rect 11057 42721 11069 42724
rect 11103 42721 11115 42755
rect 11057 42715 11115 42721
rect 21266 42712 21272 42764
rect 21324 42752 21330 42764
rect 21637 42755 21695 42761
rect 21637 42752 21649 42755
rect 21324 42724 21649 42752
rect 21324 42712 21330 42724
rect 21637 42721 21649 42724
rect 21683 42721 21695 42755
rect 21637 42715 21695 42721
rect 11330 42693 11336 42696
rect 11324 42684 11336 42693
rect 11291 42656 11336 42684
rect 11324 42647 11336 42656
rect 11330 42644 11336 42647
rect 11388 42644 11394 42696
rect 12529 42687 12587 42693
rect 12529 42653 12541 42687
rect 12575 42684 12587 42687
rect 12618 42684 12624 42696
rect 12575 42656 12624 42684
rect 12575 42653 12587 42656
rect 12529 42647 12587 42653
rect 12618 42644 12624 42656
rect 12676 42644 12682 42696
rect 12802 42644 12808 42696
rect 12860 42644 12866 42696
rect 13262 42644 13268 42696
rect 13320 42644 13326 42696
rect 13357 42687 13415 42693
rect 13357 42653 13369 42687
rect 13403 42653 13415 42687
rect 13357 42647 13415 42653
rect 13372 42616 13400 42647
rect 12728 42588 13400 42616
rect 12728 42560 12756 42588
rect 12621 42551 12679 42557
rect 12621 42517 12633 42551
rect 12667 42548 12679 42551
rect 12710 42548 12716 42560
rect 12667 42520 12716 42548
rect 12667 42517 12679 42520
rect 12621 42511 12679 42517
rect 12710 42508 12716 42520
rect 12768 42508 12774 42560
rect 12986 42508 12992 42560
rect 13044 42508 13050 42560
rect 20806 42508 20812 42560
rect 20864 42548 20870 42560
rect 21085 42551 21143 42557
rect 21085 42548 21097 42551
rect 20864 42520 21097 42548
rect 20864 42508 20870 42520
rect 21085 42517 21097 42520
rect 21131 42517 21143 42551
rect 21085 42511 21143 42517
rect 1104 42458 28888 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 28888 42458
rect 1104 42384 28888 42406
rect 12986 42168 12992 42220
rect 13044 42208 13050 42220
rect 13081 42211 13139 42217
rect 13081 42208 13093 42211
rect 13044 42180 13093 42208
rect 13044 42168 13050 42180
rect 13081 42177 13093 42180
rect 13127 42177 13139 42211
rect 13081 42171 13139 42177
rect 12529 42007 12587 42013
rect 12529 41973 12541 42007
rect 12575 42004 12587 42007
rect 12618 42004 12624 42016
rect 12575 41976 12624 42004
rect 12575 41973 12587 41976
rect 12529 41967 12587 41973
rect 12618 41964 12624 41976
rect 12676 41964 12682 42016
rect 1104 41914 28888 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 28888 41914
rect 1104 41840 28888 41862
rect 20162 41760 20168 41812
rect 20220 41760 20226 41812
rect 20257 41735 20315 41741
rect 20257 41701 20269 41735
rect 20303 41732 20315 41735
rect 20625 41735 20683 41741
rect 20625 41732 20637 41735
rect 20303 41704 20637 41732
rect 20303 41701 20315 41704
rect 20257 41695 20315 41701
rect 20625 41701 20637 41704
rect 20671 41701 20683 41735
rect 20625 41695 20683 41701
rect 17126 41556 17132 41608
rect 17184 41556 17190 41608
rect 20162 41556 20168 41608
rect 20220 41556 20226 41608
rect 20622 41556 20628 41608
rect 20680 41556 20686 41608
rect 20806 41556 20812 41608
rect 20864 41556 20870 41608
rect 22830 41556 22836 41608
rect 22888 41556 22894 41608
rect 26510 41556 26516 41608
rect 26568 41596 26574 41608
rect 26605 41599 26663 41605
rect 26605 41596 26617 41599
rect 26568 41568 26617 41596
rect 26568 41556 26574 41568
rect 26605 41565 26617 41568
rect 26651 41565 26663 41599
rect 26605 41559 26663 41565
rect 26786 41556 26792 41608
rect 26844 41556 26850 41608
rect 16666 41488 16672 41540
rect 16724 41528 16730 41540
rect 16862 41531 16920 41537
rect 16862 41528 16874 41531
rect 16724 41500 16874 41528
rect 16724 41488 16730 41500
rect 16862 41497 16874 41500
rect 16908 41497 16920 41531
rect 16862 41491 16920 41497
rect 20530 41488 20536 41540
rect 20588 41488 20594 41540
rect 23100 41531 23158 41537
rect 23100 41497 23112 41531
rect 23146 41528 23158 41531
rect 23474 41528 23480 41540
rect 23146 41500 23480 41528
rect 23146 41497 23158 41500
rect 23100 41491 23158 41497
rect 23474 41488 23480 41500
rect 23532 41488 23538 41540
rect 15749 41463 15807 41469
rect 15749 41429 15761 41463
rect 15795 41460 15807 41463
rect 17034 41460 17040 41472
rect 15795 41432 17040 41460
rect 15795 41429 15807 41432
rect 15749 41423 15807 41429
rect 17034 41420 17040 41432
rect 17092 41420 17098 41472
rect 20441 41463 20499 41469
rect 20441 41429 20453 41463
rect 20487 41460 20499 41463
rect 21082 41460 21088 41472
rect 20487 41432 21088 41460
rect 20487 41429 20499 41432
rect 20441 41423 20499 41429
rect 21082 41420 21088 41432
rect 21140 41420 21146 41472
rect 24213 41463 24271 41469
rect 24213 41429 24225 41463
rect 24259 41460 24271 41463
rect 24394 41460 24400 41472
rect 24259 41432 24400 41460
rect 24259 41429 24271 41432
rect 24213 41423 24271 41429
rect 24394 41420 24400 41432
rect 24452 41420 24458 41472
rect 26694 41420 26700 41472
rect 26752 41420 26758 41472
rect 1104 41370 28888 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 28888 41370
rect 1104 41296 28888 41318
rect 16666 41216 16672 41268
rect 16724 41216 16730 41268
rect 23474 41216 23480 41268
rect 23532 41216 23538 41268
rect 23753 41259 23811 41265
rect 23753 41225 23765 41259
rect 23799 41225 23811 41259
rect 23753 41219 23811 41225
rect 16574 41148 16580 41200
rect 16632 41188 16638 41200
rect 17221 41191 17279 41197
rect 17221 41188 17233 41191
rect 16632 41160 17233 41188
rect 16632 41148 16638 41160
rect 17221 41157 17233 41160
rect 17267 41188 17279 41191
rect 19610 41188 19616 41200
rect 17267 41160 19616 41188
rect 17267 41157 17279 41160
rect 17221 41151 17279 41157
rect 19610 41148 19616 41160
rect 19668 41188 19674 41200
rect 19668 41160 20208 41188
rect 19668 41148 19674 41160
rect 20180 41132 20208 41160
rect 16853 41123 16911 41129
rect 16853 41089 16865 41123
rect 16899 41089 16911 41123
rect 16853 41083 16911 41089
rect 17405 41123 17463 41129
rect 17405 41089 17417 41123
rect 17451 41089 17463 41123
rect 17405 41083 17463 41089
rect 17497 41123 17555 41129
rect 17497 41089 17509 41123
rect 17543 41120 17555 41123
rect 17586 41120 17592 41132
rect 17543 41092 17592 41120
rect 17543 41089 17555 41092
rect 17497 41083 17555 41089
rect 16868 40984 16896 41083
rect 17034 41012 17040 41064
rect 17092 41052 17098 41064
rect 17129 41055 17187 41061
rect 17129 41052 17141 41055
rect 17092 41024 17141 41052
rect 17092 41012 17098 41024
rect 17129 41021 17141 41024
rect 17175 41052 17187 41055
rect 17420 41052 17448 41083
rect 17586 41080 17592 41092
rect 17644 41080 17650 41132
rect 20162 41080 20168 41132
rect 20220 41120 20226 41132
rect 23382 41120 23388 41132
rect 20220 41092 23388 41120
rect 20220 41080 20226 41092
rect 23382 41080 23388 41092
rect 23440 41080 23446 41132
rect 23569 41123 23627 41129
rect 23569 41089 23581 41123
rect 23615 41120 23627 41123
rect 23768 41120 23796 41219
rect 26694 41148 26700 41200
rect 26752 41188 26758 41200
rect 27218 41191 27276 41197
rect 27218 41188 27230 41191
rect 26752 41160 27230 41188
rect 26752 41148 26758 41160
rect 27218 41157 27230 41160
rect 27264 41157 27276 41191
rect 27218 41151 27276 41157
rect 23615 41092 23796 41120
rect 23615 41089 23627 41092
rect 23569 41083 23627 41089
rect 24118 41080 24124 41132
rect 24176 41080 24182 41132
rect 26418 41080 26424 41132
rect 26476 41080 26482 41132
rect 17175 41024 17448 41052
rect 17175 41021 17187 41024
rect 17129 41015 17187 41021
rect 23198 41012 23204 41064
rect 23256 41052 23262 41064
rect 24213 41055 24271 41061
rect 24213 41052 24225 41055
rect 23256 41024 24225 41052
rect 23256 41012 23262 41024
rect 24213 41021 24225 41024
rect 24259 41021 24271 41055
rect 24213 41015 24271 41021
rect 24397 41055 24455 41061
rect 24397 41021 24409 41055
rect 24443 41052 24455 41055
rect 24578 41052 24584 41064
rect 24443 41024 24584 41052
rect 24443 41021 24455 41024
rect 24397 41015 24455 41021
rect 17221 40987 17279 40993
rect 17221 40984 17233 40987
rect 16868 40956 17233 40984
rect 17221 40953 17233 40956
rect 17267 40953 17279 40987
rect 17221 40947 17279 40953
rect 21174 40944 21180 40996
rect 21232 40984 21238 40996
rect 24412 40984 24440 41015
rect 24578 41012 24584 41024
rect 24636 41012 24642 41064
rect 26142 41012 26148 41064
rect 26200 41052 26206 41064
rect 26329 41055 26387 41061
rect 26329 41052 26341 41055
rect 26200 41024 26341 41052
rect 26200 41012 26206 41024
rect 26329 41021 26341 41024
rect 26375 41021 26387 41055
rect 26329 41015 26387 41021
rect 26970 41012 26976 41064
rect 27028 41012 27034 41064
rect 21232 40956 24440 40984
rect 21232 40944 21238 40956
rect 17037 40919 17095 40925
rect 17037 40885 17049 40919
rect 17083 40916 17095 40919
rect 17586 40916 17592 40928
rect 17083 40888 17592 40916
rect 17083 40885 17095 40888
rect 17037 40879 17095 40885
rect 17586 40876 17592 40888
rect 17644 40876 17650 40928
rect 26697 40919 26755 40925
rect 26697 40885 26709 40919
rect 26743 40916 26755 40919
rect 27154 40916 27160 40928
rect 26743 40888 27160 40916
rect 26743 40885 26755 40888
rect 26697 40879 26755 40885
rect 27154 40876 27160 40888
rect 27212 40876 27218 40928
rect 27706 40876 27712 40928
rect 27764 40916 27770 40928
rect 28353 40919 28411 40925
rect 28353 40916 28365 40919
rect 27764 40888 28365 40916
rect 27764 40876 27770 40888
rect 28353 40885 28365 40888
rect 28399 40885 28411 40919
rect 28353 40879 28411 40885
rect 1104 40826 28888 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 28888 40826
rect 1104 40752 28888 40774
rect 20441 40715 20499 40721
rect 20441 40681 20453 40715
rect 20487 40712 20499 40715
rect 20530 40712 20536 40724
rect 20487 40684 20536 40712
rect 20487 40681 20499 40684
rect 20441 40675 20499 40681
rect 20530 40672 20536 40684
rect 20588 40672 20594 40724
rect 21082 40672 21088 40724
rect 21140 40672 21146 40724
rect 23198 40672 23204 40724
rect 23256 40672 23262 40724
rect 24210 40712 24216 40724
rect 23768 40684 24216 40712
rect 20622 40604 20628 40656
rect 20680 40644 20686 40656
rect 21174 40644 21180 40656
rect 20680 40616 21180 40644
rect 20680 40604 20686 40616
rect 21174 40604 21180 40616
rect 21232 40604 21238 40656
rect 17586 40468 17592 40520
rect 17644 40508 17650 40520
rect 20640 40517 20668 40604
rect 20809 40579 20867 40585
rect 20809 40545 20821 40579
rect 20855 40576 20867 40579
rect 21082 40576 21088 40588
rect 20855 40548 21088 40576
rect 20855 40545 20867 40548
rect 20809 40539 20867 40545
rect 21082 40536 21088 40548
rect 21140 40576 21146 40588
rect 22925 40579 22983 40585
rect 21140 40548 21220 40576
rect 21140 40536 21146 40548
rect 20625 40511 20683 40517
rect 20625 40508 20637 40511
rect 17644 40480 20637 40508
rect 17644 40468 17650 40480
rect 20625 40477 20637 40480
rect 20671 40477 20683 40511
rect 20625 40471 20683 40477
rect 20901 40511 20959 40517
rect 20901 40477 20913 40511
rect 20947 40508 20959 40511
rect 20990 40508 20996 40520
rect 20947 40480 20996 40508
rect 20947 40477 20959 40480
rect 20901 40471 20959 40477
rect 20990 40468 20996 40480
rect 21048 40468 21054 40520
rect 21192 40517 21220 40548
rect 22925 40545 22937 40579
rect 22971 40576 22983 40579
rect 23474 40576 23480 40588
rect 22971 40548 23480 40576
rect 22971 40545 22983 40548
rect 22925 40539 22983 40545
rect 23474 40536 23480 40548
rect 23532 40536 23538 40588
rect 23768 40585 23796 40684
rect 24210 40672 24216 40684
rect 24268 40712 24274 40724
rect 26602 40712 26608 40724
rect 24268 40684 26608 40712
rect 24268 40672 24274 40684
rect 26602 40672 26608 40684
rect 26660 40672 26666 40724
rect 26697 40715 26755 40721
rect 26697 40681 26709 40715
rect 26743 40712 26755 40715
rect 26786 40712 26792 40724
rect 26743 40684 26792 40712
rect 26743 40681 26755 40684
rect 26697 40675 26755 40681
rect 26786 40672 26792 40684
rect 26844 40672 26850 40724
rect 23753 40579 23811 40585
rect 23753 40545 23765 40579
rect 23799 40545 23811 40579
rect 26694 40576 26700 40588
rect 23753 40539 23811 40545
rect 26436 40548 26700 40576
rect 21177 40511 21235 40517
rect 21177 40477 21189 40511
rect 21223 40477 21235 40511
rect 21177 40471 21235 40477
rect 22833 40511 22891 40517
rect 22833 40477 22845 40511
rect 22879 40508 22891 40511
rect 23661 40511 23719 40517
rect 22879 40480 23336 40508
rect 22879 40477 22891 40480
rect 22833 40471 22891 40477
rect 23308 40381 23336 40480
rect 23661 40477 23673 40511
rect 23707 40508 23719 40511
rect 24118 40508 24124 40520
rect 23707 40480 24124 40508
rect 23707 40477 23719 40480
rect 23661 40471 23719 40477
rect 24118 40468 24124 40480
rect 24176 40508 24182 40520
rect 24176 40480 24348 40508
rect 24176 40468 24182 40480
rect 24320 40384 24348 40480
rect 24394 40468 24400 40520
rect 24452 40468 24458 40520
rect 26145 40511 26203 40517
rect 26145 40477 26157 40511
rect 26191 40508 26203 40511
rect 26326 40508 26332 40520
rect 26191 40480 26332 40508
rect 26191 40477 26203 40480
rect 26145 40471 26203 40477
rect 26326 40468 26332 40480
rect 26384 40468 26390 40520
rect 26436 40517 26464 40548
rect 26694 40536 26700 40548
rect 26752 40536 26758 40588
rect 27154 40536 27160 40588
rect 27212 40536 27218 40588
rect 27338 40536 27344 40588
rect 27396 40536 27402 40588
rect 26421 40511 26479 40517
rect 26421 40477 26433 40511
rect 26467 40477 26479 40511
rect 26421 40471 26479 40477
rect 26605 40511 26663 40517
rect 26605 40477 26617 40511
rect 26651 40508 26663 40511
rect 27430 40508 27436 40520
rect 26651 40480 27436 40508
rect 26651 40477 26663 40480
rect 26605 40471 26663 40477
rect 27430 40468 27436 40480
rect 27488 40508 27494 40520
rect 27709 40511 27767 40517
rect 27709 40508 27721 40511
rect 27488 40480 27721 40508
rect 27488 40468 27494 40480
rect 27709 40477 27721 40480
rect 27755 40477 27767 40511
rect 27709 40471 27767 40477
rect 27985 40511 28043 40517
rect 27985 40477 27997 40511
rect 28031 40477 28043 40511
rect 27985 40471 28043 40477
rect 26234 40400 26240 40452
rect 26292 40440 26298 40452
rect 28000 40440 28028 40471
rect 26292 40412 28028 40440
rect 26292 40400 26298 40412
rect 23293 40375 23351 40381
rect 23293 40341 23305 40375
rect 23339 40372 23351 40375
rect 23934 40372 23940 40384
rect 23339 40344 23940 40372
rect 23339 40341 23351 40344
rect 23293 40335 23351 40341
rect 23934 40332 23940 40344
rect 23992 40332 23998 40384
rect 24302 40332 24308 40384
rect 24360 40372 24366 40384
rect 24489 40375 24547 40381
rect 24489 40372 24501 40375
rect 24360 40344 24501 40372
rect 24360 40332 24366 40344
rect 24489 40341 24501 40344
rect 24535 40341 24547 40375
rect 24489 40335 24547 40341
rect 26053 40375 26111 40381
rect 26053 40341 26065 40375
rect 26099 40372 26111 40375
rect 27065 40375 27123 40381
rect 27065 40372 27077 40375
rect 26099 40344 27077 40372
rect 26099 40341 26111 40344
rect 26053 40335 26111 40341
rect 27065 40341 27077 40344
rect 27111 40372 27123 40375
rect 27246 40372 27252 40384
rect 27111 40344 27252 40372
rect 27111 40341 27123 40344
rect 27065 40335 27123 40341
rect 27246 40332 27252 40344
rect 27304 40332 27310 40384
rect 27522 40332 27528 40384
rect 27580 40332 27586 40384
rect 27890 40332 27896 40384
rect 27948 40332 27954 40384
rect 1104 40282 28888 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 28888 40282
rect 1104 40208 28888 40230
rect 20990 40128 20996 40180
rect 21048 40168 21054 40180
rect 21091 40171 21149 40177
rect 21091 40168 21103 40171
rect 21048 40140 21103 40168
rect 21048 40128 21054 40140
rect 21091 40137 21103 40140
rect 21137 40137 21149 40171
rect 21091 40131 21149 40137
rect 23385 40171 23443 40177
rect 23385 40137 23397 40171
rect 23431 40168 23443 40171
rect 23474 40168 23480 40180
rect 23431 40140 23480 40168
rect 23431 40137 23443 40140
rect 23385 40131 23443 40137
rect 23474 40128 23480 40140
rect 23532 40128 23538 40180
rect 23753 40171 23811 40177
rect 23753 40137 23765 40171
rect 23799 40168 23811 40171
rect 26142 40168 26148 40180
rect 23799 40140 26148 40168
rect 23799 40137 23811 40140
rect 23753 40131 23811 40137
rect 26142 40128 26148 40140
rect 26200 40128 26206 40180
rect 26418 40128 26424 40180
rect 26476 40168 26482 40180
rect 26973 40171 27031 40177
rect 26973 40168 26985 40171
rect 26476 40140 26985 40168
rect 26476 40128 26482 40140
rect 26973 40137 26985 40140
rect 27019 40137 27031 40171
rect 26973 40131 27031 40137
rect 27890 40128 27896 40180
rect 27948 40128 27954 40180
rect 9582 40060 9588 40112
rect 9640 40100 9646 40112
rect 10597 40103 10655 40109
rect 10597 40100 10609 40103
rect 9640 40072 10609 40100
rect 9640 40060 9646 40072
rect 10597 40069 10609 40072
rect 10643 40069 10655 40103
rect 21177 40103 21235 40109
rect 21177 40100 21189 40103
rect 10597 40063 10655 40069
rect 20824 40072 21189 40100
rect 10612 40032 10640 40063
rect 20824 40044 20852 40072
rect 21177 40069 21189 40072
rect 21223 40069 21235 40103
rect 21177 40063 21235 40069
rect 23860 40072 24072 40100
rect 11054 40032 11060 40044
rect 10612 40004 11060 40032
rect 11054 39992 11060 40004
rect 11112 40032 11118 40044
rect 12066 40032 12072 40044
rect 11112 40004 12072 40032
rect 11112 39992 11118 40004
rect 12066 39992 12072 40004
rect 12124 39992 12130 40044
rect 12336 40035 12394 40041
rect 12336 40001 12348 40035
rect 12382 40032 12394 40035
rect 12618 40032 12624 40044
rect 12382 40004 12624 40032
rect 12382 40001 12394 40004
rect 12336 39995 12394 40001
rect 12618 39992 12624 40004
rect 12676 39992 12682 40044
rect 19797 40035 19855 40041
rect 19797 40001 19809 40035
rect 19843 40032 19855 40035
rect 19886 40032 19892 40044
rect 19843 40004 19892 40032
rect 19843 40001 19855 40004
rect 19797 39995 19855 40001
rect 19886 39992 19892 40004
rect 19944 39992 19950 40044
rect 19981 40035 20039 40041
rect 19981 40001 19993 40035
rect 20027 40032 20039 40035
rect 20070 40032 20076 40044
rect 20027 40004 20076 40032
rect 20027 40001 20039 40004
rect 19981 39995 20039 40001
rect 20070 39992 20076 40004
rect 20128 39992 20134 40044
rect 20625 40035 20683 40041
rect 20625 40001 20637 40035
rect 20671 40001 20683 40035
rect 20625 39995 20683 40001
rect 9306 39924 9312 39976
rect 9364 39924 9370 39976
rect 20162 39856 20168 39908
rect 20220 39896 20226 39908
rect 20640 39896 20668 39995
rect 20806 39992 20812 40044
rect 20864 39992 20870 40044
rect 20990 39992 20996 40044
rect 21048 39992 21054 40044
rect 21269 40035 21327 40041
rect 21269 40001 21281 40035
rect 21315 40032 21327 40035
rect 21358 40032 21364 40044
rect 21315 40004 21364 40032
rect 21315 40001 21327 40004
rect 21269 39995 21327 40001
rect 21358 39992 21364 40004
rect 21416 39992 21422 40044
rect 23106 39992 23112 40044
rect 23164 40032 23170 40044
rect 23201 40035 23259 40041
rect 23201 40032 23213 40035
rect 23164 40004 23213 40032
rect 23164 39992 23170 40004
rect 23201 40001 23213 40004
rect 23247 40001 23259 40035
rect 23201 39995 23259 40001
rect 20901 39967 20959 39973
rect 20901 39933 20913 39967
rect 20947 39933 20959 39967
rect 20901 39927 20959 39933
rect 20220 39868 20668 39896
rect 20916 39896 20944 39927
rect 21266 39896 21272 39908
rect 20916 39868 21272 39896
rect 20220 39856 20226 39868
rect 20640 39840 20668 39868
rect 21266 39856 21272 39868
rect 21324 39896 21330 39908
rect 21634 39896 21640 39908
rect 21324 39868 21640 39896
rect 21324 39856 21330 39868
rect 21634 39856 21640 39868
rect 21692 39856 21698 39908
rect 23216 39896 23244 39995
rect 23290 39992 23296 40044
rect 23348 40032 23354 40044
rect 23860 40032 23888 40072
rect 23348 40004 23888 40032
rect 23348 39992 23354 40004
rect 23934 39992 23940 40044
rect 23992 39992 23998 40044
rect 24044 40032 24072 40072
rect 27430 40060 27436 40112
rect 27488 40060 27494 40112
rect 27706 40060 27712 40112
rect 27764 40060 27770 40112
rect 24121 40035 24179 40041
rect 24121 40032 24133 40035
rect 24044 40004 24133 40032
rect 24121 40001 24133 40004
rect 24167 40001 24179 40035
rect 24121 39995 24179 40001
rect 24394 39992 24400 40044
rect 24452 39992 24458 40044
rect 24670 39992 24676 40044
rect 24728 40032 24734 40044
rect 26234 40032 26240 40044
rect 24728 40004 26240 40032
rect 24728 39992 24734 40004
rect 26234 39992 26240 40004
rect 26292 39992 26298 40044
rect 26694 39992 26700 40044
rect 26752 40032 26758 40044
rect 27525 40035 27583 40041
rect 27525 40032 27537 40035
rect 26752 40004 27537 40032
rect 26752 39992 26758 40004
rect 27525 40001 27537 40004
rect 27571 40001 27583 40035
rect 27525 39995 27583 40001
rect 23658 39924 23664 39976
rect 23716 39924 23722 39976
rect 24029 39967 24087 39973
rect 24029 39933 24041 39967
rect 24075 39933 24087 39967
rect 24029 39927 24087 39933
rect 24213 39967 24271 39973
rect 24213 39933 24225 39967
rect 24259 39964 24271 39967
rect 24857 39967 24915 39973
rect 24857 39964 24869 39967
rect 24259 39936 24869 39964
rect 24259 39933 24271 39936
rect 24213 39927 24271 39933
rect 24857 39933 24869 39936
rect 24903 39933 24915 39967
rect 24857 39927 24915 39933
rect 24044 39896 24072 39927
rect 23216 39868 24072 39896
rect 27157 39899 27215 39905
rect 27157 39865 27169 39899
rect 27203 39896 27215 39899
rect 27890 39896 27896 39908
rect 27203 39868 27896 39896
rect 27203 39865 27215 39868
rect 27157 39859 27215 39865
rect 27890 39856 27896 39868
rect 27948 39856 27954 39908
rect 8478 39788 8484 39840
rect 8536 39828 8542 39840
rect 8757 39831 8815 39837
rect 8757 39828 8769 39831
rect 8536 39800 8769 39828
rect 8536 39788 8542 39800
rect 8757 39797 8769 39800
rect 8803 39797 8815 39831
rect 8757 39791 8815 39797
rect 13446 39788 13452 39840
rect 13504 39788 13510 39840
rect 19794 39788 19800 39840
rect 19852 39828 19858 39840
rect 19981 39831 20039 39837
rect 19981 39828 19993 39831
rect 19852 39800 19993 39828
rect 19852 39788 19858 39800
rect 19981 39797 19993 39800
rect 20027 39797 20039 39831
rect 19981 39791 20039 39797
rect 20438 39788 20444 39840
rect 20496 39788 20502 39840
rect 20622 39788 20628 39840
rect 20680 39828 20686 39840
rect 21358 39828 21364 39840
rect 20680 39800 21364 39828
rect 20680 39788 20686 39800
rect 21358 39788 21364 39800
rect 21416 39788 21422 39840
rect 24026 39788 24032 39840
rect 24084 39828 24090 39840
rect 24489 39831 24547 39837
rect 24489 39828 24501 39831
rect 24084 39800 24501 39828
rect 24084 39788 24090 39800
rect 24489 39797 24501 39800
rect 24535 39797 24547 39831
rect 24489 39791 24547 39797
rect 1104 39738 28888 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 28888 39738
rect 1104 39664 28888 39686
rect 10965 39627 11023 39633
rect 10965 39593 10977 39627
rect 11011 39624 11023 39627
rect 11054 39624 11060 39636
rect 11011 39596 11060 39624
rect 11011 39593 11023 39596
rect 10965 39587 11023 39593
rect 11054 39584 11060 39596
rect 11112 39584 11118 39636
rect 17402 39584 17408 39636
rect 17460 39624 17466 39636
rect 17586 39624 17592 39636
rect 17460 39596 17592 39624
rect 17460 39584 17466 39596
rect 17586 39584 17592 39596
rect 17644 39584 17650 39636
rect 18049 39627 18107 39633
rect 18049 39593 18061 39627
rect 18095 39624 18107 39627
rect 18322 39624 18328 39636
rect 18095 39596 18328 39624
rect 18095 39593 18107 39596
rect 18049 39587 18107 39593
rect 18322 39584 18328 39596
rect 18380 39624 18386 39636
rect 20162 39624 20168 39636
rect 18380 39596 20168 39624
rect 18380 39584 18386 39596
rect 20162 39584 20168 39596
rect 20220 39584 20226 39636
rect 20257 39627 20315 39633
rect 20257 39593 20269 39627
rect 20303 39624 20315 39627
rect 20990 39624 20996 39636
rect 20303 39596 20996 39624
rect 20303 39593 20315 39596
rect 20257 39587 20315 39593
rect 20272 39556 20300 39587
rect 20990 39584 20996 39596
rect 21048 39584 21054 39636
rect 21082 39584 21088 39636
rect 21140 39584 21146 39636
rect 21266 39584 21272 39636
rect 21324 39624 21330 39636
rect 23566 39624 23572 39636
rect 21324 39596 23572 39624
rect 21324 39584 21330 39596
rect 23566 39584 23572 39596
rect 23624 39584 23630 39636
rect 23658 39584 23664 39636
rect 23716 39624 23722 39636
rect 24121 39627 24179 39633
rect 24121 39624 24133 39627
rect 23716 39596 24133 39624
rect 23716 39584 23722 39596
rect 24121 39593 24133 39596
rect 24167 39624 24179 39627
rect 24167 39596 24900 39624
rect 24167 39593 24179 39596
rect 24121 39587 24179 39593
rect 19628 39528 20300 39556
rect 12066 39448 12072 39500
rect 12124 39488 12130 39500
rect 12529 39491 12587 39497
rect 12529 39488 12541 39491
rect 12124 39460 12541 39488
rect 12124 39448 12130 39460
rect 12529 39457 12541 39460
rect 12575 39457 12587 39491
rect 12529 39451 12587 39457
rect 16758 39448 16764 39500
rect 16816 39448 16822 39500
rect 17034 39488 17040 39500
rect 16868 39460 17040 39488
rect 8478 39380 8484 39432
rect 8536 39380 8542 39432
rect 8573 39423 8631 39429
rect 8573 39389 8585 39423
rect 8619 39389 8631 39423
rect 8573 39383 8631 39389
rect 8588 39284 8616 39383
rect 8938 39380 8944 39432
rect 8996 39420 9002 39432
rect 9582 39420 9588 39432
rect 8996 39392 9588 39420
rect 8996 39380 9002 39392
rect 9582 39380 9588 39392
rect 9640 39380 9646 39432
rect 12434 39420 12440 39432
rect 9692 39392 12440 39420
rect 8757 39355 8815 39361
rect 8757 39321 8769 39355
rect 8803 39352 8815 39355
rect 9186 39355 9244 39361
rect 9186 39352 9198 39355
rect 8803 39324 9198 39352
rect 8803 39321 8815 39324
rect 8757 39315 8815 39321
rect 9186 39321 9198 39324
rect 9232 39321 9244 39355
rect 9186 39315 9244 39321
rect 9692 39296 9720 39392
rect 12434 39380 12440 39392
rect 12492 39420 12498 39432
rect 13354 39420 13360 39432
rect 12492 39392 13360 39420
rect 12492 39380 12498 39392
rect 13354 39380 13360 39392
rect 13412 39380 13418 39432
rect 16868 39429 16896 39460
rect 17034 39448 17040 39460
rect 17092 39488 17098 39500
rect 17092 39460 18276 39488
rect 17092 39448 17098 39460
rect 18248 39429 18276 39460
rect 19628 39429 19656 39528
rect 19904 39460 20208 39488
rect 19904 39432 19932 39460
rect 16853 39423 16911 39429
rect 16853 39389 16865 39423
rect 16899 39389 16911 39423
rect 17865 39423 17923 39429
rect 17865 39420 17877 39423
rect 16853 39383 16911 39389
rect 17604 39392 17877 39420
rect 12250 39312 12256 39364
rect 12308 39312 12314 39364
rect 12796 39355 12854 39361
rect 12796 39321 12808 39355
rect 12842 39352 12854 39355
rect 13170 39352 13176 39364
rect 12842 39324 13176 39352
rect 12842 39321 12854 39324
rect 12796 39315 12854 39321
rect 13170 39312 13176 39324
rect 13228 39312 13234 39364
rect 16206 39312 16212 39364
rect 16264 39352 16270 39364
rect 17604 39352 17632 39392
rect 17865 39389 17877 39392
rect 17911 39389 17923 39423
rect 17865 39383 17923 39389
rect 18233 39423 18291 39429
rect 18233 39389 18245 39423
rect 18279 39389 18291 39423
rect 18233 39383 18291 39389
rect 19613 39423 19671 39429
rect 19613 39389 19625 39423
rect 19659 39389 19671 39423
rect 19613 39383 19671 39389
rect 16264 39324 17632 39352
rect 17681 39355 17739 39361
rect 16264 39312 16270 39324
rect 17681 39321 17693 39355
rect 17727 39352 17739 39355
rect 17770 39352 17776 39364
rect 17727 39324 17776 39352
rect 17727 39321 17739 39324
rect 17681 39315 17739 39321
rect 17770 39312 17776 39324
rect 17828 39312 17834 39364
rect 17880 39352 17908 39383
rect 19794 39380 19800 39432
rect 19852 39380 19858 39432
rect 19886 39380 19892 39432
rect 19944 39380 19950 39432
rect 20070 39380 20076 39432
rect 20128 39380 20134 39432
rect 20180 39420 20208 39460
rect 20438 39448 20444 39500
rect 20496 39448 20502 39500
rect 20717 39491 20775 39497
rect 20717 39457 20729 39491
rect 20763 39488 20775 39491
rect 21100 39488 21128 39584
rect 24670 39556 24676 39568
rect 20763 39460 21128 39488
rect 21192 39528 21404 39556
rect 20763 39457 20775 39460
rect 20717 39451 20775 39457
rect 20533 39423 20591 39429
rect 20533 39420 20545 39423
rect 20180 39392 20545 39420
rect 20533 39389 20545 39392
rect 20579 39389 20591 39423
rect 20533 39383 20591 39389
rect 20625 39423 20683 39429
rect 20625 39389 20637 39423
rect 20671 39389 20683 39423
rect 20625 39383 20683 39389
rect 20088 39352 20116 39380
rect 20640 39352 20668 39383
rect 21192 39352 21220 39528
rect 21266 39448 21272 39500
rect 21324 39448 21330 39500
rect 21376 39488 21404 39528
rect 22066 39528 24676 39556
rect 22066 39488 22094 39528
rect 24670 39516 24676 39528
rect 24728 39516 24734 39568
rect 24765 39491 24823 39497
rect 21376 39460 22094 39488
rect 23676 39460 24256 39488
rect 21358 39380 21364 39432
rect 21416 39380 21422 39432
rect 21634 39380 21640 39432
rect 21692 39380 21698 39432
rect 17880 39324 19564 39352
rect 20088 39324 20668 39352
rect 20732 39324 21220 39352
rect 21376 39352 21404 39380
rect 21729 39355 21787 39361
rect 21729 39352 21741 39355
rect 21376 39324 21741 39352
rect 9674 39284 9680 39296
rect 8588 39256 9680 39284
rect 9674 39244 9680 39256
rect 9732 39244 9738 39296
rect 10318 39244 10324 39296
rect 10376 39244 10382 39296
rect 13909 39287 13967 39293
rect 13909 39253 13921 39287
rect 13955 39284 13967 39287
rect 14550 39284 14556 39296
rect 13955 39256 14556 39284
rect 13955 39253 13967 39256
rect 13909 39247 13967 39253
rect 14550 39244 14556 39256
rect 14608 39244 14614 39296
rect 17218 39244 17224 39296
rect 17276 39244 17282 39296
rect 18325 39287 18383 39293
rect 18325 39253 18337 39287
rect 18371 39284 18383 39287
rect 18506 39284 18512 39296
rect 18371 39256 18512 39284
rect 18371 39253 18383 39256
rect 18325 39247 18383 39253
rect 18506 39244 18512 39256
rect 18564 39244 18570 39296
rect 19426 39244 19432 39296
rect 19484 39244 19490 39296
rect 19536 39284 19564 39324
rect 20732 39284 20760 39324
rect 21729 39321 21741 39324
rect 21775 39321 21787 39355
rect 21729 39315 21787 39321
rect 23566 39312 23572 39364
rect 23624 39352 23630 39364
rect 23676 39352 23704 39460
rect 24228 39432 24256 39460
rect 24765 39457 24777 39491
rect 24811 39488 24823 39491
rect 24872 39488 24900 39596
rect 24811 39460 24900 39488
rect 24811 39457 24823 39460
rect 24765 39451 24823 39457
rect 23753 39423 23811 39429
rect 23753 39389 23765 39423
rect 23799 39420 23811 39423
rect 24026 39420 24032 39432
rect 23799 39392 24032 39420
rect 23799 39389 23811 39392
rect 23753 39383 23811 39389
rect 24026 39380 24032 39392
rect 24084 39380 24090 39432
rect 24210 39380 24216 39432
rect 24268 39380 24274 39432
rect 24581 39423 24639 39429
rect 24581 39389 24593 39423
rect 24627 39389 24639 39423
rect 24581 39383 24639 39389
rect 23624 39324 23704 39352
rect 23937 39355 23995 39361
rect 23624 39312 23630 39324
rect 23937 39321 23949 39355
rect 23983 39352 23995 39355
rect 24596 39352 24624 39383
rect 23983 39324 24624 39352
rect 23983 39321 23995 39324
rect 23937 39315 23995 39321
rect 19536 39256 20760 39284
rect 20901 39287 20959 39293
rect 20901 39253 20913 39287
rect 20947 39284 20959 39287
rect 23106 39284 23112 39296
rect 20947 39256 23112 39284
rect 20947 39253 20959 39256
rect 20901 39247 20959 39253
rect 23106 39244 23112 39256
rect 23164 39244 23170 39296
rect 23290 39244 23296 39296
rect 23348 39284 23354 39296
rect 24397 39287 24455 39293
rect 24397 39284 24409 39287
rect 23348 39256 24409 39284
rect 23348 39244 23354 39256
rect 24397 39253 24409 39256
rect 24443 39253 24455 39287
rect 24397 39247 24455 39253
rect 1104 39194 28888 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 28888 39194
rect 1104 39120 28888 39142
rect 9033 39083 9091 39089
rect 9033 39049 9045 39083
rect 9079 39080 9091 39083
rect 9306 39080 9312 39092
rect 9079 39052 9312 39080
rect 9079 39049 9091 39052
rect 9033 39043 9091 39049
rect 9306 39040 9312 39052
rect 9364 39040 9370 39092
rect 13170 39040 13176 39092
rect 13228 39040 13234 39092
rect 16206 39040 16212 39092
rect 16264 39040 16270 39092
rect 16850 39080 16856 39092
rect 16500 39052 16856 39080
rect 8938 39012 8944 39024
rect 7668 38984 8944 39012
rect 7668 38953 7696 38984
rect 8938 38972 8944 38984
rect 8996 38972 9002 39024
rect 7926 38953 7932 38956
rect 7653 38947 7711 38953
rect 7653 38913 7665 38947
rect 7699 38913 7711 38947
rect 7653 38907 7711 38913
rect 7920 38907 7932 38953
rect 7926 38904 7932 38907
rect 7984 38904 7990 38956
rect 9582 38904 9588 38956
rect 9640 38904 9646 38956
rect 9858 38953 9864 38956
rect 9852 38907 9864 38953
rect 9858 38904 9864 38907
rect 9916 38904 9922 38956
rect 13354 38904 13360 38956
rect 13412 38904 13418 38956
rect 13446 38904 13452 38956
rect 13504 38904 13510 38956
rect 14550 38904 14556 38956
rect 14608 38904 14614 38956
rect 14737 38947 14795 38953
rect 14737 38913 14749 38947
rect 14783 38913 14795 38947
rect 14737 38907 14795 38913
rect 14274 38836 14280 38888
rect 14332 38876 14338 38888
rect 14752 38876 14780 38907
rect 16022 38904 16028 38956
rect 16080 38904 16086 38956
rect 16206 38904 16212 38956
rect 16264 38904 16270 38956
rect 16500 38953 16528 39052
rect 16850 39040 16856 39052
rect 16908 39040 16914 39092
rect 18877 39083 18935 39089
rect 18877 39049 18889 39083
rect 18923 39080 18935 39083
rect 18923 39052 19288 39080
rect 18923 39049 18935 39052
rect 18877 39043 18935 39049
rect 17126 39012 17132 39024
rect 16684 38984 17132 39012
rect 16684 38953 16712 38984
rect 17126 38972 17132 38984
rect 17184 39012 17190 39024
rect 17184 38984 19104 39012
rect 17184 38972 17190 38984
rect 16301 38947 16359 38953
rect 16301 38913 16313 38947
rect 16347 38913 16359 38947
rect 16301 38907 16359 38913
rect 16485 38947 16543 38953
rect 16485 38913 16497 38947
rect 16531 38913 16543 38947
rect 16485 38907 16543 38913
rect 16669 38947 16727 38953
rect 16669 38913 16681 38947
rect 16715 38913 16727 38947
rect 16925 38947 16983 38953
rect 16925 38944 16937 38947
rect 16669 38907 16727 38913
rect 16776 38916 16937 38944
rect 14332 38848 14780 38876
rect 14332 38836 14338 38848
rect 10594 38700 10600 38752
rect 10652 38740 10658 38752
rect 10965 38743 11023 38749
rect 10965 38740 10977 38743
rect 10652 38712 10977 38740
rect 10652 38700 10658 38712
rect 10965 38709 10977 38712
rect 11011 38709 11023 38743
rect 10965 38703 11023 38709
rect 14645 38743 14703 38749
rect 14645 38709 14657 38743
rect 14691 38740 14703 38743
rect 15378 38740 15384 38752
rect 14691 38712 15384 38740
rect 14691 38709 14703 38712
rect 14645 38703 14703 38709
rect 15378 38700 15384 38712
rect 15436 38700 15442 38752
rect 16316 38740 16344 38907
rect 16393 38879 16451 38885
rect 16393 38845 16405 38879
rect 16439 38876 16451 38879
rect 16776 38876 16804 38916
rect 16925 38913 16937 38916
rect 16971 38913 16983 38947
rect 16925 38907 16983 38913
rect 18322 38904 18328 38956
rect 18380 38904 18386 38956
rect 18598 38904 18604 38956
rect 18656 38904 18662 38956
rect 16439 38848 16804 38876
rect 18509 38879 18567 38885
rect 16439 38845 16451 38848
rect 16393 38839 16451 38845
rect 18509 38845 18521 38879
rect 18555 38845 18567 38879
rect 18509 38839 18567 38845
rect 18049 38811 18107 38817
rect 18049 38777 18061 38811
rect 18095 38808 18107 38811
rect 18230 38808 18236 38820
rect 18095 38780 18236 38808
rect 18095 38777 18107 38780
rect 18049 38771 18107 38777
rect 18230 38768 18236 38780
rect 18288 38808 18294 38820
rect 18524 38808 18552 38839
rect 18874 38836 18880 38888
rect 18932 38836 18938 38888
rect 19076 38885 19104 38984
rect 19260 38944 19288 39052
rect 19426 39040 19432 39092
rect 19484 39080 19490 39092
rect 20993 39083 21051 39089
rect 20993 39080 21005 39083
rect 19484 39052 21005 39080
rect 19484 39040 19490 39052
rect 20993 39049 21005 39052
rect 21039 39049 21051 39083
rect 20993 39043 21051 39049
rect 19328 39015 19386 39021
rect 19328 38981 19340 39015
rect 19374 39012 19386 39015
rect 19518 39012 19524 39024
rect 19374 38984 19524 39012
rect 19374 38981 19386 38984
rect 19328 38975 19386 38981
rect 19518 38972 19524 38984
rect 19576 38972 19582 39024
rect 19886 38944 19892 38956
rect 19260 38916 19892 38944
rect 19886 38904 19892 38916
rect 19944 38904 19950 38956
rect 20254 38904 20260 38956
rect 20312 38944 20318 38956
rect 20901 38947 20959 38953
rect 20901 38944 20913 38947
rect 20312 38916 20913 38944
rect 20312 38904 20318 38916
rect 20901 38913 20913 38916
rect 20947 38913 20959 38947
rect 20901 38907 20959 38913
rect 23201 38947 23259 38953
rect 23201 38913 23213 38947
rect 23247 38944 23259 38947
rect 23290 38944 23296 38956
rect 23247 38916 23296 38944
rect 23247 38913 23259 38916
rect 23201 38907 23259 38913
rect 23290 38904 23296 38916
rect 23348 38904 23354 38956
rect 19061 38879 19119 38885
rect 19061 38845 19073 38879
rect 19107 38845 19119 38879
rect 19061 38839 19119 38845
rect 18288 38780 18552 38808
rect 18288 38768 18294 38780
rect 16574 38740 16580 38752
rect 16316 38712 16580 38740
rect 16574 38700 16580 38712
rect 16632 38700 16638 38752
rect 16666 38700 16672 38752
rect 16724 38740 16730 38752
rect 17770 38740 17776 38752
rect 16724 38712 17776 38740
rect 16724 38700 16730 38712
rect 17770 38700 17776 38712
rect 17828 38700 17834 38752
rect 18138 38700 18144 38752
rect 18196 38700 18202 38752
rect 18690 38700 18696 38752
rect 18748 38700 18754 38752
rect 19076 38740 19104 38839
rect 21174 38836 21180 38888
rect 21232 38836 21238 38888
rect 23106 38836 23112 38888
rect 23164 38836 23170 38888
rect 20438 38768 20444 38820
rect 20496 38808 20502 38820
rect 20806 38808 20812 38820
rect 20496 38780 20812 38808
rect 20496 38768 20502 38780
rect 20806 38768 20812 38780
rect 20864 38768 20870 38820
rect 23566 38768 23572 38820
rect 23624 38768 23630 38820
rect 19334 38740 19340 38752
rect 19076 38712 19340 38740
rect 19334 38700 19340 38712
rect 19392 38700 19398 38752
rect 20530 38700 20536 38752
rect 20588 38700 20594 38752
rect 1104 38650 28888 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 28888 38650
rect 1104 38576 28888 38598
rect 7926 38496 7932 38548
rect 7984 38536 7990 38548
rect 8113 38539 8171 38545
rect 8113 38536 8125 38539
rect 7984 38508 8125 38536
rect 7984 38496 7990 38508
rect 8113 38505 8125 38508
rect 8159 38505 8171 38539
rect 8113 38499 8171 38505
rect 9858 38496 9864 38548
rect 9916 38496 9922 38548
rect 14274 38496 14280 38548
rect 14332 38496 14338 38548
rect 15657 38539 15715 38545
rect 15657 38505 15669 38539
rect 15703 38536 15715 38539
rect 16666 38536 16672 38548
rect 15703 38508 16672 38536
rect 15703 38505 15715 38508
rect 15657 38499 15715 38505
rect 16666 38496 16672 38508
rect 16724 38496 16730 38548
rect 16758 38496 16764 38548
rect 16816 38496 16822 38548
rect 16850 38496 16856 38548
rect 16908 38496 16914 38548
rect 19518 38496 19524 38548
rect 19576 38496 19582 38548
rect 20070 38496 20076 38548
rect 20128 38496 20134 38548
rect 26878 38496 26884 38548
rect 26936 38536 26942 38548
rect 27338 38536 27344 38548
rect 26936 38508 27344 38536
rect 26936 38496 26942 38508
rect 27338 38496 27344 38508
rect 27396 38496 27402 38548
rect 13909 38471 13967 38477
rect 13909 38437 13921 38471
rect 13955 38468 13967 38471
rect 14829 38471 14887 38477
rect 13955 38440 14780 38468
rect 13955 38437 13967 38440
rect 13909 38431 13967 38437
rect 9493 38403 9551 38409
rect 9493 38369 9505 38403
rect 9539 38400 9551 38403
rect 10689 38403 10747 38409
rect 10689 38400 10701 38403
rect 9539 38372 10701 38400
rect 9539 38369 9551 38372
rect 9493 38363 9551 38369
rect 10689 38369 10701 38372
rect 10735 38369 10747 38403
rect 10689 38363 10747 38369
rect 13446 38360 13452 38412
rect 13504 38360 13510 38412
rect 14752 38400 14780 38440
rect 14829 38437 14841 38471
rect 14875 38468 14887 38471
rect 16022 38468 16028 38480
rect 14875 38440 16028 38468
rect 14875 38437 14887 38440
rect 14829 38431 14887 38437
rect 16022 38428 16028 38440
rect 16080 38428 16086 38480
rect 18138 38468 18144 38480
rect 16684 38440 18144 38468
rect 14752 38372 15700 38400
rect 8294 38292 8300 38344
rect 8352 38292 8358 38344
rect 8481 38335 8539 38341
rect 8481 38301 8493 38335
rect 8527 38332 8539 38335
rect 8570 38332 8576 38344
rect 8527 38304 8576 38332
rect 8527 38301 8539 38304
rect 8481 38295 8539 38301
rect 8570 38292 8576 38304
rect 8628 38292 8634 38344
rect 9674 38292 9680 38344
rect 9732 38292 9738 38344
rect 10594 38292 10600 38344
rect 10652 38292 10658 38344
rect 11241 38335 11299 38341
rect 11241 38301 11253 38335
rect 11287 38301 11299 38335
rect 11241 38295 11299 38301
rect 10318 38224 10324 38276
rect 10376 38264 10382 38276
rect 11256 38264 11284 38295
rect 12526 38292 12532 38344
rect 12584 38332 12590 38344
rect 13541 38335 13599 38341
rect 13541 38332 13553 38335
rect 12584 38304 13553 38332
rect 12584 38292 12590 38304
rect 13541 38301 13553 38304
rect 13587 38332 13599 38335
rect 13722 38332 13728 38344
rect 13587 38304 13728 38332
rect 13587 38301 13599 38304
rect 13541 38295 13599 38301
rect 13722 38292 13728 38304
rect 13780 38332 13786 38344
rect 14185 38335 14243 38341
rect 14185 38332 14197 38335
rect 13780 38304 14197 38332
rect 13780 38292 13786 38304
rect 14185 38301 14197 38304
rect 14231 38301 14243 38335
rect 14185 38295 14243 38301
rect 14550 38292 14556 38344
rect 14608 38292 14614 38344
rect 14642 38292 14648 38344
rect 14700 38292 14706 38344
rect 15378 38292 15384 38344
rect 15436 38292 15442 38344
rect 15672 38341 15700 38372
rect 15657 38335 15715 38341
rect 15657 38301 15669 38335
rect 15703 38301 15715 38335
rect 15657 38295 15715 38301
rect 16577 38335 16635 38341
rect 16577 38301 16589 38335
rect 16623 38332 16635 38335
rect 16684 38332 16712 38440
rect 18138 38428 18144 38440
rect 18196 38428 18202 38480
rect 20530 38468 20536 38480
rect 19628 38440 20536 38468
rect 17218 38360 17224 38412
rect 17276 38400 17282 38412
rect 17313 38403 17371 38409
rect 17313 38400 17325 38403
rect 17276 38372 17325 38400
rect 17276 38360 17282 38372
rect 17313 38369 17325 38372
rect 17359 38369 17371 38403
rect 17313 38363 17371 38369
rect 17402 38360 17408 38412
rect 17460 38360 17466 38412
rect 18690 38400 18696 38412
rect 17512 38372 18696 38400
rect 16623 38304 16712 38332
rect 16761 38335 16819 38341
rect 16623 38301 16635 38304
rect 16577 38295 16635 38301
rect 16761 38301 16773 38335
rect 16807 38332 16819 38335
rect 16942 38332 16948 38344
rect 16807 38304 16948 38332
rect 16807 38301 16819 38304
rect 16761 38295 16819 38301
rect 16942 38292 16948 38304
rect 17000 38332 17006 38344
rect 17512 38332 17540 38372
rect 18690 38360 18696 38372
rect 18748 38360 18754 38412
rect 17000 38304 17540 38332
rect 17000 38292 17006 38304
rect 17678 38292 17684 38344
rect 17736 38292 17742 38344
rect 17957 38335 18015 38341
rect 17957 38301 17969 38335
rect 18003 38301 18015 38335
rect 17957 38295 18015 38301
rect 10376 38236 11284 38264
rect 14568 38264 14596 38292
rect 14921 38267 14979 38273
rect 14921 38264 14933 38267
rect 14568 38236 14933 38264
rect 10376 38224 10382 38236
rect 14921 38233 14933 38236
rect 14967 38233 14979 38267
rect 14921 38227 14979 38233
rect 15105 38267 15163 38273
rect 15105 38233 15117 38267
rect 15151 38233 15163 38267
rect 17773 38267 17831 38273
rect 17773 38264 17785 38267
rect 15105 38227 15163 38233
rect 16776 38236 17785 38264
rect 9953 38199 10011 38205
rect 9953 38165 9965 38199
rect 9999 38196 10011 38199
rect 10134 38196 10140 38208
rect 9999 38168 10140 38196
rect 9999 38165 10011 38168
rect 9953 38159 10011 38165
rect 10134 38156 10140 38168
rect 10192 38156 10198 38208
rect 14274 38156 14280 38208
rect 14332 38196 14338 38208
rect 15120 38196 15148 38227
rect 14332 38168 15148 38196
rect 15289 38199 15347 38205
rect 14332 38156 14338 38168
rect 15289 38165 15301 38199
rect 15335 38196 15347 38199
rect 15473 38199 15531 38205
rect 15473 38196 15485 38199
rect 15335 38168 15485 38196
rect 15335 38165 15347 38168
rect 15289 38159 15347 38165
rect 15473 38165 15485 38168
rect 15519 38165 15531 38199
rect 15473 38159 15531 38165
rect 16206 38156 16212 38208
rect 16264 38196 16270 38208
rect 16482 38196 16488 38208
rect 16264 38168 16488 38196
rect 16264 38156 16270 38168
rect 16482 38156 16488 38168
rect 16540 38196 16546 38208
rect 16776 38196 16804 38236
rect 17773 38233 17785 38236
rect 17819 38233 17831 38267
rect 17773 38227 17831 38233
rect 16540 38168 16804 38196
rect 17221 38199 17279 38205
rect 16540 38156 16546 38168
rect 17221 38165 17233 38199
rect 17267 38196 17279 38199
rect 17972 38196 18000 38295
rect 18230 38292 18236 38344
rect 18288 38292 18294 38344
rect 19337 38335 19395 38341
rect 19337 38301 19349 38335
rect 19383 38301 19395 38335
rect 19337 38295 19395 38301
rect 19521 38335 19579 38341
rect 19521 38301 19533 38335
rect 19567 38332 19579 38335
rect 19628 38332 19656 38440
rect 20530 38428 20536 38440
rect 20588 38428 20594 38480
rect 19889 38403 19947 38409
rect 19889 38369 19901 38403
rect 19935 38400 19947 38403
rect 20622 38400 20628 38412
rect 19935 38372 20628 38400
rect 19935 38369 19947 38372
rect 19889 38363 19947 38369
rect 20622 38360 20628 38372
rect 20680 38360 20686 38412
rect 27154 38360 27160 38412
rect 27212 38360 27218 38412
rect 19567 38304 19656 38332
rect 19797 38335 19855 38341
rect 19567 38301 19579 38304
rect 19521 38295 19579 38301
rect 19797 38301 19809 38335
rect 19843 38332 19855 38335
rect 19843 38304 20300 38332
rect 19843 38301 19855 38304
rect 19797 38295 19855 38301
rect 18141 38267 18199 38273
rect 18141 38233 18153 38267
rect 18187 38264 18199 38267
rect 18874 38264 18880 38276
rect 18187 38236 18880 38264
rect 18187 38233 18199 38236
rect 18141 38227 18199 38233
rect 18874 38224 18880 38236
rect 18932 38224 18938 38276
rect 19352 38264 19380 38295
rect 19610 38264 19616 38276
rect 19352 38236 19616 38264
rect 19610 38224 19616 38236
rect 19668 38224 19674 38276
rect 20272 38208 20300 38304
rect 20438 38292 20444 38344
rect 20496 38332 20502 38344
rect 20533 38335 20591 38341
rect 20533 38332 20545 38335
rect 20496 38304 20545 38332
rect 20496 38292 20502 38304
rect 20533 38301 20545 38304
rect 20579 38301 20591 38335
rect 20533 38295 20591 38301
rect 27065 38335 27123 38341
rect 27065 38301 27077 38335
rect 27111 38332 27123 38335
rect 27522 38332 27528 38344
rect 27111 38304 27528 38332
rect 27111 38301 27123 38304
rect 27065 38295 27123 38301
rect 27522 38292 27528 38304
rect 27580 38292 27586 38344
rect 18322 38196 18328 38208
rect 17267 38168 18328 38196
rect 17267 38165 17279 38168
rect 17221 38159 17279 38165
rect 18322 38156 18328 38168
rect 18380 38156 18386 38208
rect 20254 38156 20260 38208
rect 20312 38196 20318 38208
rect 20441 38199 20499 38205
rect 20441 38196 20453 38199
rect 20312 38168 20453 38196
rect 20312 38156 20318 38168
rect 20441 38165 20453 38168
rect 20487 38165 20499 38199
rect 20441 38159 20499 38165
rect 26697 38199 26755 38205
rect 26697 38165 26709 38199
rect 26743 38196 26755 38199
rect 27062 38196 27068 38208
rect 26743 38168 27068 38196
rect 26743 38165 26755 38168
rect 26697 38159 26755 38165
rect 27062 38156 27068 38168
rect 27120 38156 27126 38208
rect 1104 38106 28888 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 28888 38106
rect 1104 38032 28888 38054
rect 8570 37952 8576 38004
rect 8628 37952 8634 38004
rect 9769 37995 9827 38001
rect 9769 37961 9781 37995
rect 9815 37992 9827 37995
rect 10594 37992 10600 38004
rect 9815 37964 10600 37992
rect 9815 37961 9827 37964
rect 9769 37955 9827 37961
rect 10594 37952 10600 37964
rect 10652 37952 10658 38004
rect 16022 37952 16028 38004
rect 16080 37992 16086 38004
rect 17113 37995 17171 38001
rect 17113 37992 17125 37995
rect 16080 37964 17125 37992
rect 16080 37952 16086 37964
rect 17113 37961 17125 37964
rect 17159 37992 17171 37995
rect 17678 37992 17684 38004
rect 17159 37964 17684 37992
rect 17159 37961 17171 37964
rect 17113 37955 17171 37961
rect 17678 37952 17684 37964
rect 17736 37952 17742 38004
rect 17770 37952 17776 38004
rect 17828 37992 17834 38004
rect 17828 37964 18460 37992
rect 17828 37952 17834 37964
rect 9306 37884 9312 37936
rect 9364 37924 9370 37936
rect 9493 37927 9551 37933
rect 9493 37924 9505 37927
rect 9364 37896 9505 37924
rect 9364 37884 9370 37896
rect 9493 37893 9505 37896
rect 9539 37893 9551 37927
rect 9493 37887 9551 37893
rect 9861 37927 9919 37933
rect 9861 37893 9873 37927
rect 9907 37924 9919 37927
rect 10318 37924 10324 37936
rect 9907 37896 10324 37924
rect 9907 37893 9919 37896
rect 9861 37887 9919 37893
rect 10318 37884 10324 37896
rect 10376 37884 10382 37936
rect 12434 37884 12440 37936
rect 12492 37924 12498 37936
rect 12618 37924 12624 37936
rect 12492 37896 12624 37924
rect 12492 37884 12498 37896
rect 12618 37884 12624 37896
rect 12676 37884 12682 37936
rect 14550 37924 14556 37936
rect 14200 37896 14556 37924
rect 9217 37859 9275 37865
rect 9217 37825 9229 37859
rect 9263 37856 9275 37859
rect 9674 37856 9680 37868
rect 9263 37828 9680 37856
rect 9263 37825 9275 37828
rect 9217 37819 9275 37825
rect 9674 37816 9680 37828
rect 9732 37816 9738 37868
rect 12253 37859 12311 37865
rect 12253 37856 12265 37859
rect 10336 37828 12265 37856
rect 8478 37748 8484 37800
rect 8536 37788 8542 37800
rect 10336 37788 10364 37828
rect 12253 37825 12265 37828
rect 12299 37856 12311 37859
rect 12805 37859 12863 37865
rect 12805 37856 12817 37859
rect 12299 37828 12817 37856
rect 12299 37825 12311 37828
rect 12253 37819 12311 37825
rect 12805 37825 12817 37828
rect 12851 37856 12863 37859
rect 13262 37856 13268 37868
rect 12851 37828 13268 37856
rect 12851 37825 12863 37828
rect 12805 37819 12863 37825
rect 13262 37816 13268 37828
rect 13320 37816 13326 37868
rect 13722 37816 13728 37868
rect 13780 37856 13786 37868
rect 14200 37865 14228 37896
rect 14550 37884 14556 37896
rect 14608 37884 14614 37936
rect 17313 37927 17371 37933
rect 17313 37893 17325 37927
rect 17359 37924 17371 37927
rect 18322 37924 18328 37936
rect 17359 37896 18328 37924
rect 17359 37893 17371 37896
rect 17313 37887 17371 37893
rect 18322 37884 18328 37896
rect 18380 37884 18386 37936
rect 18432 37924 18460 37964
rect 19610 37952 19616 38004
rect 19668 37992 19674 38004
rect 20530 37992 20536 38004
rect 19668 37964 20536 37992
rect 19668 37952 19674 37964
rect 20530 37952 20536 37964
rect 20588 37952 20594 38004
rect 23566 37952 23572 38004
rect 23624 37992 23630 38004
rect 23753 37995 23811 38001
rect 23753 37992 23765 37995
rect 23624 37964 23765 37992
rect 23624 37952 23630 37964
rect 23753 37961 23765 37964
rect 23799 37961 23811 37995
rect 23753 37955 23811 37961
rect 26973 37995 27031 38001
rect 26973 37961 26985 37995
rect 27019 37992 27031 37995
rect 27154 37992 27160 38004
rect 27019 37964 27160 37992
rect 27019 37961 27031 37964
rect 26973 37955 27031 37961
rect 27154 37952 27160 37964
rect 27212 37952 27218 38004
rect 18432 37896 27200 37924
rect 27172 37868 27200 37896
rect 14093 37859 14151 37865
rect 14093 37856 14105 37859
rect 13780 37828 14105 37856
rect 13780 37816 13786 37828
rect 14093 37825 14105 37828
rect 14139 37825 14151 37859
rect 14093 37819 14151 37825
rect 14185 37859 14243 37865
rect 14185 37825 14197 37859
rect 14231 37825 14243 37859
rect 14185 37819 14243 37825
rect 14274 37816 14280 37868
rect 14332 37816 14338 37868
rect 14369 37859 14427 37865
rect 14369 37825 14381 37859
rect 14415 37856 14427 37859
rect 14642 37856 14648 37868
rect 14415 37828 14648 37856
rect 14415 37825 14427 37828
rect 14369 37819 14427 37825
rect 8536 37760 10364 37788
rect 8536 37748 8542 37760
rect 11146 37748 11152 37800
rect 11204 37748 11210 37800
rect 12529 37791 12587 37797
rect 12529 37757 12541 37791
rect 12575 37788 12587 37791
rect 12710 37788 12716 37800
rect 12575 37760 12716 37788
rect 12575 37757 12587 37760
rect 12529 37751 12587 37757
rect 12710 37748 12716 37760
rect 12768 37748 12774 37800
rect 13446 37748 13452 37800
rect 13504 37788 13510 37800
rect 14384 37788 14412 37819
rect 14642 37816 14648 37828
rect 14700 37816 14706 37868
rect 23658 37816 23664 37868
rect 23716 37816 23722 37868
rect 27154 37816 27160 37868
rect 27212 37816 27218 37868
rect 27338 37816 27344 37868
rect 27396 37816 27402 37868
rect 13504 37760 14412 37788
rect 14553 37791 14611 37797
rect 13504 37748 13510 37760
rect 14553 37757 14565 37791
rect 14599 37788 14611 37791
rect 16482 37788 16488 37800
rect 14599 37760 16488 37788
rect 14599 37757 14611 37760
rect 14553 37751 14611 37757
rect 16482 37748 16488 37760
rect 16540 37788 16546 37800
rect 23937 37791 23995 37797
rect 16540 37748 16574 37788
rect 23937 37757 23949 37791
rect 23983 37757 23995 37791
rect 23937 37751 23995 37757
rect 16546 37720 16574 37748
rect 23952 37720 23980 37751
rect 26234 37748 26240 37800
rect 26292 37788 26298 37800
rect 27249 37791 27307 37797
rect 27249 37788 27261 37791
rect 26292 37760 27261 37788
rect 26292 37748 26298 37760
rect 27249 37757 27261 37760
rect 27295 37757 27307 37791
rect 27249 37751 27307 37757
rect 24578 37720 24584 37732
rect 16546 37692 17172 37720
rect 23952 37692 24584 37720
rect 9766 37612 9772 37664
rect 9824 37652 9830 37664
rect 10045 37655 10103 37661
rect 10045 37652 10057 37655
rect 9824 37624 10057 37652
rect 9824 37612 9830 37624
rect 10045 37621 10057 37624
rect 10091 37621 10103 37655
rect 10045 37615 10103 37621
rect 10502 37612 10508 37664
rect 10560 37652 10566 37664
rect 10597 37655 10655 37661
rect 10597 37652 10609 37655
rect 10560 37624 10609 37652
rect 10560 37612 10566 37624
rect 10597 37621 10609 37624
rect 10643 37621 10655 37655
rect 10597 37615 10655 37621
rect 16942 37612 16948 37664
rect 17000 37612 17006 37664
rect 17144 37661 17172 37692
rect 24578 37680 24584 37692
rect 24636 37720 24642 37732
rect 26878 37720 26884 37732
rect 24636 37692 26884 37720
rect 24636 37680 24642 37692
rect 26878 37680 26884 37692
rect 26936 37680 26942 37732
rect 17129 37655 17187 37661
rect 17129 37621 17141 37655
rect 17175 37621 17187 37655
rect 17129 37615 17187 37621
rect 23290 37612 23296 37664
rect 23348 37612 23354 37664
rect 1104 37562 28888 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 28888 37562
rect 1104 37488 28888 37510
rect 8294 37408 8300 37460
rect 8352 37448 8358 37460
rect 8941 37451 8999 37457
rect 8941 37448 8953 37451
rect 8352 37420 8953 37448
rect 8352 37408 8358 37420
rect 8941 37417 8953 37420
rect 8987 37417 8999 37451
rect 8941 37411 8999 37417
rect 10134 37408 10140 37460
rect 10192 37408 10198 37460
rect 23750 37408 23756 37460
rect 23808 37448 23814 37460
rect 24489 37451 24547 37457
rect 24489 37448 24501 37451
rect 23808 37420 24501 37448
rect 23808 37408 23814 37420
rect 24489 37417 24501 37420
rect 24535 37417 24547 37451
rect 24489 37411 24547 37417
rect 8665 37383 8723 37389
rect 8665 37349 8677 37383
rect 8711 37380 8723 37383
rect 9674 37380 9680 37392
rect 8711 37352 9680 37380
rect 8711 37349 8723 37352
rect 8665 37343 8723 37349
rect 9674 37340 9680 37352
rect 9732 37340 9738 37392
rect 26789 37383 26847 37389
rect 26789 37349 26801 37383
rect 26835 37380 26847 37383
rect 27157 37383 27215 37389
rect 27157 37380 27169 37383
rect 26835 37352 27169 37380
rect 26835 37349 26847 37352
rect 26789 37343 26847 37349
rect 27157 37349 27169 37352
rect 27203 37349 27215 37383
rect 27157 37343 27215 37349
rect 9306 37312 9312 37324
rect 8956 37284 9312 37312
rect 7285 37247 7343 37253
rect 7285 37213 7297 37247
rect 7331 37244 7343 37247
rect 8386 37244 8392 37256
rect 7331 37216 8392 37244
rect 7331 37213 7343 37216
rect 7285 37207 7343 37213
rect 8386 37204 8392 37216
rect 8444 37204 8450 37256
rect 8956 37253 8984 37284
rect 9306 37272 9312 37284
rect 9364 37272 9370 37324
rect 10318 37272 10324 37324
rect 10376 37272 10382 37324
rect 8941 37247 8999 37253
rect 8941 37213 8953 37247
rect 8987 37213 8999 37247
rect 8941 37207 8999 37213
rect 9125 37247 9183 37253
rect 9125 37213 9137 37247
rect 9171 37213 9183 37247
rect 9125 37207 9183 37213
rect 7552 37179 7610 37185
rect 7552 37145 7564 37179
rect 7598 37176 7610 37179
rect 8018 37176 8024 37188
rect 7598 37148 8024 37176
rect 7598 37145 7610 37148
rect 7552 37139 7610 37145
rect 8018 37136 8024 37148
rect 8076 37136 8082 37188
rect 9140 37176 9168 37207
rect 9214 37204 9220 37256
rect 9272 37204 9278 37256
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 10413 37247 10471 37253
rect 10413 37244 10425 37247
rect 9732 37216 10425 37244
rect 9732 37204 9738 37216
rect 10413 37213 10425 37216
rect 10459 37213 10471 37247
rect 10413 37207 10471 37213
rect 10689 37247 10747 37253
rect 10689 37213 10701 37247
rect 10735 37244 10747 37247
rect 12161 37247 12219 37253
rect 12161 37244 12173 37247
rect 10735 37216 12173 37244
rect 10735 37213 10747 37216
rect 10689 37207 10747 37213
rect 11072 37188 11100 37216
rect 12161 37213 12173 37216
rect 12207 37213 12219 37247
rect 12161 37207 12219 37213
rect 22830 37204 22836 37256
rect 22888 37244 22894 37256
rect 22888 37216 24348 37244
rect 22888 37204 22894 37216
rect 9306 37176 9312 37188
rect 9140 37148 9312 37176
rect 9306 37136 9312 37148
rect 9364 37136 9370 37188
rect 10962 37185 10968 37188
rect 10137 37179 10195 37185
rect 10137 37145 10149 37179
rect 10183 37145 10195 37179
rect 10137 37139 10195 37145
rect 10956 37139 10968 37185
rect 9401 37111 9459 37117
rect 9401 37077 9413 37111
rect 9447 37108 9459 37111
rect 10152 37108 10180 37139
rect 10962 37136 10968 37139
rect 11020 37136 11026 37188
rect 11054 37136 11060 37188
rect 11112 37136 11118 37188
rect 12434 37185 12440 37188
rect 12428 37139 12440 37185
rect 12434 37136 12440 37139
rect 12492 37136 12498 37188
rect 23100 37179 23158 37185
rect 23100 37145 23112 37179
rect 23146 37176 23158 37179
rect 23198 37176 23204 37188
rect 23146 37148 23204 37176
rect 23146 37145 23158 37148
rect 23100 37139 23158 37145
rect 23198 37136 23204 37148
rect 23256 37136 23262 37188
rect 24320 37176 24348 37216
rect 24394 37204 24400 37256
rect 24452 37204 24458 37256
rect 26510 37204 26516 37256
rect 26568 37244 26574 37256
rect 26697 37247 26755 37253
rect 26697 37244 26709 37247
rect 26568 37216 26709 37244
rect 26568 37204 26574 37216
rect 26697 37213 26709 37216
rect 26743 37213 26755 37247
rect 26697 37207 26755 37213
rect 26878 37204 26884 37256
rect 26936 37204 26942 37256
rect 27062 37204 27068 37256
rect 27120 37204 27126 37256
rect 27154 37204 27160 37256
rect 27212 37204 27218 37256
rect 27341 37247 27399 37253
rect 27341 37213 27353 37247
rect 27387 37244 27399 37247
rect 27893 37247 27951 37253
rect 27893 37244 27905 37247
rect 27387 37216 27905 37244
rect 27387 37213 27399 37216
rect 27341 37207 27399 37213
rect 27893 37213 27905 37216
rect 27939 37213 27951 37247
rect 27893 37207 27951 37213
rect 28442 37204 28448 37256
rect 28500 37204 28506 37256
rect 24320 37148 24624 37176
rect 9447 37080 10180 37108
rect 10597 37111 10655 37117
rect 9447 37077 9459 37080
rect 9401 37071 9459 37077
rect 10597 37077 10609 37111
rect 10643 37108 10655 37111
rect 11146 37108 11152 37120
rect 10643 37080 11152 37108
rect 10643 37077 10655 37080
rect 10597 37071 10655 37077
rect 11146 37068 11152 37080
rect 11204 37068 11210 37120
rect 12069 37111 12127 37117
rect 12069 37077 12081 37111
rect 12115 37108 12127 37111
rect 12526 37108 12532 37120
rect 12115 37080 12532 37108
rect 12115 37077 12127 37080
rect 12069 37071 12127 37077
rect 12526 37068 12532 37080
rect 12584 37068 12590 37120
rect 13541 37111 13599 37117
rect 13541 37077 13553 37111
rect 13587 37108 13599 37111
rect 14274 37108 14280 37120
rect 13587 37080 14280 37108
rect 13587 37077 13599 37080
rect 13541 37071 13599 37077
rect 14274 37068 14280 37080
rect 14332 37068 14338 37120
rect 24026 37068 24032 37120
rect 24084 37108 24090 37120
rect 24213 37111 24271 37117
rect 24213 37108 24225 37111
rect 24084 37080 24225 37108
rect 24084 37068 24090 37080
rect 24213 37077 24225 37080
rect 24259 37108 24271 37111
rect 24394 37108 24400 37120
rect 24259 37080 24400 37108
rect 24259 37077 24271 37080
rect 24213 37071 24271 37077
rect 24394 37068 24400 37080
rect 24452 37068 24458 37120
rect 24596 37108 24624 37148
rect 26602 37136 26608 37188
rect 26660 37136 26666 37188
rect 26878 37108 26884 37120
rect 24596 37080 26884 37108
rect 26878 37068 26884 37080
rect 26936 37068 26942 37120
rect 1104 37018 28888 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 28888 37018
rect 1104 36944 28888 36966
rect 8018 36864 8024 36916
rect 8076 36864 8082 36916
rect 9769 36907 9827 36913
rect 9769 36904 9781 36907
rect 9416 36876 9781 36904
rect 8205 36771 8263 36777
rect 8205 36737 8217 36771
rect 8251 36768 8263 36771
rect 8478 36768 8484 36780
rect 8251 36740 8484 36768
rect 8251 36737 8263 36740
rect 8205 36731 8263 36737
rect 8478 36728 8484 36740
rect 8536 36728 8542 36780
rect 8389 36703 8447 36709
rect 8389 36669 8401 36703
rect 8435 36700 8447 36703
rect 8849 36703 8907 36709
rect 8849 36700 8861 36703
rect 8435 36672 8861 36700
rect 8435 36669 8447 36672
rect 8389 36663 8447 36669
rect 8849 36669 8861 36672
rect 8895 36669 8907 36703
rect 8849 36663 8907 36669
rect 9306 36660 9312 36712
rect 9364 36700 9370 36712
rect 9416 36709 9444 36876
rect 9769 36873 9781 36876
rect 9815 36873 9827 36907
rect 9769 36867 9827 36873
rect 10873 36907 10931 36913
rect 10873 36873 10885 36907
rect 10919 36904 10931 36907
rect 10962 36904 10968 36916
rect 10919 36876 10968 36904
rect 10919 36873 10931 36876
rect 10873 36867 10931 36873
rect 10962 36864 10968 36876
rect 11020 36864 11026 36916
rect 12253 36907 12311 36913
rect 12253 36873 12265 36907
rect 12299 36904 12311 36907
rect 12434 36904 12440 36916
rect 12299 36876 12440 36904
rect 12299 36873 12311 36876
rect 12253 36867 12311 36873
rect 10502 36796 10508 36848
rect 10560 36796 10566 36848
rect 10597 36839 10655 36845
rect 10597 36805 10609 36839
rect 10643 36836 10655 36839
rect 11790 36836 11796 36848
rect 10643 36808 11796 36836
rect 10643 36805 10655 36808
rect 10597 36799 10655 36805
rect 11790 36796 11796 36808
rect 11848 36796 11854 36848
rect 9585 36771 9643 36777
rect 9585 36737 9597 36771
rect 9631 36768 9643 36771
rect 9766 36768 9772 36780
rect 9631 36740 9772 36768
rect 9631 36737 9643 36740
rect 9585 36731 9643 36737
rect 9766 36728 9772 36740
rect 9824 36728 9830 36780
rect 10045 36771 10103 36777
rect 10045 36737 10057 36771
rect 10091 36768 10103 36771
rect 10321 36771 10379 36777
rect 10321 36768 10333 36771
rect 10091 36740 10333 36768
rect 10091 36737 10103 36740
rect 10045 36731 10103 36737
rect 9401 36703 9459 36709
rect 9401 36700 9413 36703
rect 9364 36672 9413 36700
rect 9364 36660 9370 36672
rect 9401 36669 9413 36672
rect 9447 36669 9459 36703
rect 9401 36663 9459 36669
rect 9674 36660 9680 36712
rect 9732 36660 9738 36712
rect 9953 36703 10011 36709
rect 9953 36669 9965 36703
rect 9999 36669 10011 36703
rect 9953 36663 10011 36669
rect 8294 36592 8300 36644
rect 8352 36632 8358 36644
rect 9968 36632 9996 36663
rect 8352 36604 9996 36632
rect 10152 36632 10180 36740
rect 10321 36737 10333 36740
rect 10367 36737 10379 36771
rect 10321 36731 10379 36737
rect 10689 36771 10747 36777
rect 10689 36737 10701 36771
rect 10735 36737 10747 36771
rect 10689 36731 10747 36737
rect 10229 36703 10287 36709
rect 10229 36669 10241 36703
rect 10275 36700 10287 36703
rect 10704 36700 10732 36731
rect 10275 36672 10732 36700
rect 10275 36669 10287 36672
rect 10229 36663 10287 36669
rect 12268 36632 12296 36867
rect 12434 36864 12440 36876
rect 12492 36864 12498 36916
rect 23198 36864 23204 36916
rect 23256 36864 23262 36916
rect 26697 36907 26755 36913
rect 26697 36873 26709 36907
rect 26743 36904 26755 36907
rect 27338 36904 27344 36916
rect 26743 36876 27344 36904
rect 26743 36873 26755 36876
rect 26697 36867 26755 36873
rect 27338 36864 27344 36876
rect 27396 36864 27402 36916
rect 12618 36836 12624 36848
rect 12452 36808 12624 36836
rect 12452 36777 12480 36808
rect 12618 36796 12624 36808
rect 12676 36796 12682 36848
rect 23382 36836 23388 36848
rect 23124 36808 23388 36836
rect 12437 36771 12495 36777
rect 12437 36737 12449 36771
rect 12483 36737 12495 36771
rect 12437 36731 12495 36737
rect 12526 36728 12532 36780
rect 12584 36728 12590 36780
rect 19334 36728 19340 36780
rect 19392 36768 19398 36780
rect 20901 36771 20959 36777
rect 20901 36768 20913 36771
rect 19392 36740 20913 36768
rect 19392 36728 19398 36740
rect 20901 36737 20913 36740
rect 20947 36768 20959 36771
rect 22830 36768 22836 36780
rect 20947 36740 22836 36768
rect 20947 36737 20959 36740
rect 20901 36731 20959 36737
rect 22830 36728 22836 36740
rect 22888 36728 22894 36780
rect 23124 36777 23152 36808
rect 23382 36796 23388 36808
rect 23440 36796 23446 36848
rect 26602 36796 26608 36848
rect 26660 36836 26666 36848
rect 27218 36839 27276 36845
rect 27218 36836 27230 36839
rect 26660 36808 27230 36836
rect 26660 36796 26666 36808
rect 27218 36805 27230 36808
rect 27264 36805 27276 36839
rect 27218 36799 27276 36805
rect 23109 36771 23167 36777
rect 23109 36737 23121 36771
rect 23155 36737 23167 36771
rect 23109 36731 23167 36737
rect 23290 36728 23296 36780
rect 23348 36728 23354 36780
rect 26789 36771 26847 36777
rect 26789 36737 26801 36771
rect 26835 36737 26847 36771
rect 26789 36731 26847 36737
rect 10152 36604 12296 36632
rect 8352 36592 8358 36604
rect 26804 36564 26832 36731
rect 26970 36728 26976 36780
rect 27028 36728 27034 36780
rect 28353 36567 28411 36573
rect 28353 36564 28365 36567
rect 26804 36536 28365 36564
rect 28353 36533 28365 36536
rect 28399 36564 28411 36567
rect 28442 36564 28448 36576
rect 28399 36536 28448 36564
rect 28399 36533 28411 36536
rect 28353 36527 28411 36533
rect 28442 36524 28448 36536
rect 28500 36524 28506 36576
rect 1104 36474 28888 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 28888 36474
rect 1104 36400 28888 36422
rect 9214 36184 9220 36236
rect 9272 36224 9278 36236
rect 9490 36224 9496 36236
rect 9272 36196 9496 36224
rect 9272 36184 9278 36196
rect 9490 36184 9496 36196
rect 9548 36184 9554 36236
rect 22189 36227 22247 36233
rect 22189 36193 22201 36227
rect 22235 36224 22247 36227
rect 22830 36224 22836 36236
rect 22235 36196 22836 36224
rect 22235 36193 22247 36196
rect 22189 36187 22247 36193
rect 22830 36184 22836 36196
rect 22888 36184 22894 36236
rect 12250 36048 12256 36100
rect 12308 36088 12314 36100
rect 19886 36088 19892 36100
rect 12308 36060 19892 36088
rect 12308 36048 12314 36060
rect 19886 36048 19892 36060
rect 19944 36088 19950 36100
rect 20441 36091 20499 36097
rect 20441 36088 20453 36091
rect 19944 36060 20453 36088
rect 19944 36048 19950 36060
rect 20441 36057 20453 36060
rect 20487 36057 20499 36091
rect 20441 36051 20499 36057
rect 8938 35980 8944 36032
rect 8996 35980 9002 36032
rect 1104 35930 28888 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 28888 35930
rect 1104 35856 28888 35878
rect 6914 35816 6920 35828
rect 6564 35788 6920 35816
rect 6564 35689 6592 35788
rect 6914 35776 6920 35788
rect 6972 35816 6978 35828
rect 6972 35788 9076 35816
rect 6972 35776 6978 35788
rect 8386 35748 8392 35760
rect 6840 35720 8392 35748
rect 6840 35689 6868 35720
rect 8386 35708 8392 35720
rect 8444 35708 8450 35760
rect 6549 35683 6607 35689
rect 6549 35649 6561 35683
rect 6595 35649 6607 35683
rect 6549 35643 6607 35649
rect 6825 35683 6883 35689
rect 6825 35649 6837 35683
rect 6871 35649 6883 35683
rect 7081 35683 7139 35689
rect 7081 35680 7093 35683
rect 6825 35643 6883 35649
rect 6932 35652 7093 35680
rect 6362 35572 6368 35624
rect 6420 35572 6426 35624
rect 6733 35615 6791 35621
rect 6733 35581 6745 35615
rect 6779 35612 6791 35615
rect 6932 35612 6960 35652
rect 7081 35649 7093 35652
rect 7127 35649 7139 35683
rect 7081 35643 7139 35649
rect 8938 35640 8944 35692
rect 8996 35640 9002 35692
rect 9048 35689 9076 35788
rect 9306 35776 9312 35828
rect 9364 35776 9370 35828
rect 9217 35751 9275 35757
rect 9217 35717 9229 35751
rect 9263 35748 9275 35751
rect 9674 35748 9680 35760
rect 9263 35720 9680 35748
rect 9263 35717 9275 35720
rect 9217 35711 9275 35717
rect 9674 35708 9680 35720
rect 9732 35708 9738 35760
rect 12066 35748 12072 35760
rect 9784 35720 12072 35748
rect 9033 35683 9091 35689
rect 9033 35649 9045 35683
rect 9079 35680 9091 35683
rect 9784 35680 9812 35720
rect 12066 35708 12072 35720
rect 12124 35708 12130 35760
rect 18598 35708 18604 35760
rect 18656 35748 18662 35760
rect 19521 35751 19579 35757
rect 19521 35748 19533 35751
rect 18656 35720 19533 35748
rect 18656 35708 18662 35720
rect 19521 35717 19533 35720
rect 19567 35717 19579 35751
rect 19521 35711 19579 35717
rect 9079 35652 9812 35680
rect 10433 35683 10491 35689
rect 9079 35649 9091 35652
rect 9033 35643 9091 35649
rect 10433 35649 10445 35683
rect 10479 35680 10491 35683
rect 11882 35680 11888 35692
rect 10479 35652 11888 35680
rect 10479 35649 10491 35652
rect 10433 35643 10491 35649
rect 11882 35640 11888 35652
rect 11940 35640 11946 35692
rect 18874 35640 18880 35692
rect 18932 35680 18938 35692
rect 19429 35683 19487 35689
rect 19429 35680 19441 35683
rect 18932 35652 19441 35680
rect 18932 35640 18938 35652
rect 19429 35649 19441 35652
rect 19475 35649 19487 35683
rect 19429 35643 19487 35649
rect 19705 35683 19763 35689
rect 19705 35649 19717 35683
rect 19751 35680 19763 35683
rect 20346 35680 20352 35692
rect 19751 35652 20352 35680
rect 19751 35649 19763 35652
rect 19705 35643 19763 35649
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 28258 35640 28264 35692
rect 28316 35640 28322 35692
rect 6779 35584 6960 35612
rect 6779 35581 6791 35584
rect 6733 35575 6791 35581
rect 10686 35572 10692 35624
rect 10744 35572 10750 35624
rect 26786 35572 26792 35624
rect 26844 35612 26850 35624
rect 26973 35615 27031 35621
rect 26973 35612 26985 35615
rect 26844 35584 26985 35612
rect 26844 35572 26850 35584
rect 26973 35581 26985 35584
rect 27019 35581 27031 35615
rect 26973 35575 27031 35581
rect 8205 35547 8263 35553
rect 8205 35513 8217 35547
rect 8251 35544 8263 35547
rect 9490 35544 9496 35556
rect 8251 35516 9496 35544
rect 8251 35513 8263 35516
rect 8205 35507 8263 35513
rect 9490 35504 9496 35516
rect 9548 35504 9554 35556
rect 19705 35479 19763 35485
rect 19705 35445 19717 35479
rect 19751 35476 19763 35479
rect 20714 35476 20720 35488
rect 19751 35448 20720 35476
rect 19751 35445 19763 35448
rect 19705 35439 19763 35445
rect 20714 35436 20720 35448
rect 20772 35436 20778 35488
rect 27614 35436 27620 35488
rect 27672 35436 27678 35488
rect 28442 35436 28448 35488
rect 28500 35436 28506 35488
rect 1104 35386 28888 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 28888 35386
rect 1104 35312 28888 35334
rect 6362 35232 6368 35284
rect 6420 35232 6426 35284
rect 11790 35232 11796 35284
rect 11848 35232 11854 35284
rect 11882 35232 11888 35284
rect 11940 35232 11946 35284
rect 28258 35232 28264 35284
rect 28316 35232 28322 35284
rect 7006 35096 7012 35148
rect 7064 35136 7070 35148
rect 8294 35136 8300 35148
rect 7064 35108 8300 35136
rect 7064 35096 7070 35108
rect 8294 35096 8300 35108
rect 8352 35096 8358 35148
rect 11808 35136 11836 35232
rect 18874 35164 18880 35216
rect 18932 35204 18938 35216
rect 18932 35176 19840 35204
rect 18932 35164 18938 35176
rect 12253 35139 12311 35145
rect 12253 35136 12265 35139
rect 11808 35108 12265 35136
rect 12253 35105 12265 35108
rect 12299 35105 12311 35139
rect 12253 35099 12311 35105
rect 19518 35096 19524 35148
rect 19576 35096 19582 35148
rect 11146 35028 11152 35080
rect 11204 35028 11210 35080
rect 12066 35028 12072 35080
rect 12124 35028 12130 35080
rect 19426 35028 19432 35080
rect 19484 35028 19490 35080
rect 19812 35077 19840 35176
rect 19705 35071 19763 35077
rect 19705 35037 19717 35071
rect 19751 35037 19763 35071
rect 19705 35031 19763 35037
rect 19797 35071 19855 35077
rect 19797 35037 19809 35071
rect 19843 35037 19855 35071
rect 19797 35031 19855 35037
rect 19981 35071 20039 35077
rect 19981 35037 19993 35071
rect 20027 35068 20039 35071
rect 20073 35071 20131 35077
rect 20073 35068 20085 35071
rect 20027 35040 20085 35068
rect 20027 35037 20039 35040
rect 19981 35031 20039 35037
rect 20073 35037 20085 35040
rect 20119 35037 20131 35071
rect 20073 35031 20131 35037
rect 20349 35071 20407 35077
rect 20349 35037 20361 35071
rect 20395 35068 20407 35071
rect 20806 35068 20812 35080
rect 20395 35040 20812 35068
rect 20395 35037 20407 35040
rect 20349 35031 20407 35037
rect 8386 34960 8392 35012
rect 8444 34960 8450 35012
rect 9309 35003 9367 35009
rect 9309 34969 9321 35003
rect 9355 35000 9367 35003
rect 12158 35000 12164 35012
rect 9355 34972 12164 35000
rect 9355 34969 9367 34972
rect 9309 34963 9367 34969
rect 12158 34960 12164 34972
rect 12216 34960 12222 35012
rect 18322 34960 18328 35012
rect 18380 35000 18386 35012
rect 19720 35000 19748 35031
rect 20806 35028 20812 35040
rect 20864 35028 20870 35080
rect 20898 35028 20904 35080
rect 20956 35028 20962 35080
rect 26881 35071 26939 35077
rect 26881 35037 26893 35071
rect 26927 35068 26939 35071
rect 26970 35068 26976 35080
rect 26927 35040 26976 35068
rect 26927 35037 26939 35040
rect 26881 35031 26939 35037
rect 26970 35028 26976 35040
rect 27028 35028 27034 35080
rect 27148 35071 27206 35077
rect 27148 35037 27160 35071
rect 27194 35068 27206 35071
rect 27614 35068 27620 35080
rect 27194 35040 27620 35068
rect 27194 35037 27206 35040
rect 27148 35031 27206 35037
rect 27614 35028 27620 35040
rect 27672 35028 27678 35080
rect 18380 34972 19748 35000
rect 20533 35003 20591 35009
rect 18380 34960 18386 34972
rect 20533 34969 20545 35003
rect 20579 35000 20591 35003
rect 22002 35000 22008 35012
rect 20579 34972 22008 35000
rect 20579 34969 20591 34972
rect 20533 34963 20591 34969
rect 22002 34960 22008 34972
rect 22060 34960 22066 35012
rect 8404 34932 8432 34960
rect 8846 34932 8852 34944
rect 8404 34904 8852 34932
rect 8846 34892 8852 34904
rect 8904 34932 8910 34944
rect 10597 34935 10655 34941
rect 10597 34932 10609 34935
rect 8904 34904 10609 34932
rect 8904 34892 8910 34904
rect 10597 34901 10609 34904
rect 10643 34932 10655 34935
rect 10686 34932 10692 34944
rect 10643 34904 10692 34932
rect 10643 34901 10655 34904
rect 10597 34895 10655 34901
rect 10686 34892 10692 34904
rect 10744 34892 10750 34944
rect 19334 34892 19340 34944
rect 19392 34932 19398 34944
rect 20165 34935 20223 34941
rect 20165 34932 20177 34935
rect 19392 34904 20177 34932
rect 19392 34892 19398 34904
rect 20165 34901 20177 34904
rect 20211 34901 20223 34935
rect 20165 34895 20223 34901
rect 20622 34892 20628 34944
rect 20680 34932 20686 34944
rect 20717 34935 20775 34941
rect 20717 34932 20729 34935
rect 20680 34904 20729 34932
rect 20680 34892 20686 34904
rect 20717 34901 20729 34904
rect 20763 34932 20775 34935
rect 20990 34932 20996 34944
rect 20763 34904 20996 34932
rect 20763 34901 20775 34904
rect 20717 34895 20775 34901
rect 20990 34892 20996 34904
rect 21048 34892 21054 34944
rect 1104 34842 28888 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 28888 34842
rect 1104 34768 28888 34790
rect 6181 34731 6239 34737
rect 6181 34697 6193 34731
rect 6227 34728 6239 34731
rect 7006 34728 7012 34740
rect 6227 34700 7012 34728
rect 6227 34697 6239 34700
rect 6181 34691 6239 34697
rect 7006 34688 7012 34700
rect 7064 34688 7070 34740
rect 10689 34731 10747 34737
rect 10689 34697 10701 34731
rect 10735 34728 10747 34731
rect 11146 34728 11152 34740
rect 10735 34700 11152 34728
rect 10735 34697 10747 34700
rect 10689 34691 10747 34697
rect 11146 34688 11152 34700
rect 11204 34688 11210 34740
rect 20346 34688 20352 34740
rect 20404 34688 20410 34740
rect 20806 34688 20812 34740
rect 20864 34728 20870 34740
rect 21637 34731 21695 34737
rect 21637 34728 21649 34731
rect 20864 34700 21649 34728
rect 20864 34688 20870 34700
rect 21637 34697 21649 34700
rect 21683 34697 21695 34731
rect 21637 34691 21695 34697
rect 24121 34731 24179 34737
rect 24121 34697 24133 34731
rect 24167 34728 24179 34731
rect 25222 34728 25228 34740
rect 24167 34700 25228 34728
rect 24167 34697 24179 34700
rect 24121 34691 24179 34697
rect 25222 34688 25228 34700
rect 25280 34688 25286 34740
rect 26421 34731 26479 34737
rect 26421 34697 26433 34731
rect 26467 34728 26479 34731
rect 27338 34728 27344 34740
rect 26467 34700 27344 34728
rect 26467 34697 26479 34700
rect 26421 34691 26479 34697
rect 27338 34688 27344 34700
rect 27396 34688 27402 34740
rect 9576 34663 9634 34669
rect 4816 34632 6914 34660
rect 4816 34601 4844 34632
rect 4801 34595 4859 34601
rect 4801 34561 4813 34595
rect 4847 34561 4859 34595
rect 5057 34595 5115 34601
rect 5057 34592 5069 34595
rect 4801 34555 4859 34561
rect 4908 34564 5069 34592
rect 4614 34484 4620 34536
rect 4672 34524 4678 34536
rect 4908 34524 4936 34564
rect 5057 34561 5069 34564
rect 5103 34561 5115 34595
rect 5057 34555 5115 34561
rect 4672 34496 4936 34524
rect 6886 34524 6914 34632
rect 9576 34629 9588 34663
rect 9622 34660 9634 34663
rect 9674 34660 9680 34672
rect 9622 34632 9680 34660
rect 9622 34629 9634 34632
rect 9576 34623 9634 34629
rect 9674 34620 9680 34632
rect 9732 34620 9738 34672
rect 18322 34620 18328 34672
rect 18380 34660 18386 34672
rect 18380 34632 18828 34660
rect 18380 34620 18386 34632
rect 16206 34552 16212 34604
rect 16264 34601 16270 34604
rect 16264 34555 16276 34601
rect 16264 34552 16270 34555
rect 18506 34552 18512 34604
rect 18564 34552 18570 34604
rect 18598 34552 18604 34604
rect 18656 34552 18662 34604
rect 18800 34601 18828 34632
rect 21358 34620 21364 34672
rect 21416 34660 21422 34672
rect 21416 34632 22324 34660
rect 21416 34620 21422 34632
rect 18785 34595 18843 34601
rect 18785 34561 18797 34595
rect 18831 34561 18843 34595
rect 18785 34555 18843 34561
rect 18874 34552 18880 34604
rect 18932 34552 18938 34604
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 20254 34592 20260 34604
rect 19484 34564 20260 34592
rect 19484 34552 19490 34564
rect 20254 34552 20260 34564
rect 20312 34592 20318 34604
rect 21085 34595 21143 34601
rect 21085 34592 21097 34595
rect 20312 34564 21097 34592
rect 20312 34552 20318 34564
rect 21085 34561 21097 34564
rect 21131 34561 21143 34595
rect 21085 34555 21143 34561
rect 21269 34595 21327 34601
rect 21269 34561 21281 34595
rect 21315 34561 21327 34595
rect 21269 34555 21327 34561
rect 21453 34595 21511 34601
rect 21453 34561 21465 34595
rect 21499 34561 21511 34595
rect 21453 34555 21511 34561
rect 8846 34524 8852 34536
rect 6886 34496 8852 34524
rect 4672 34484 4678 34496
rect 8846 34484 8852 34496
rect 8904 34524 8910 34536
rect 9309 34527 9367 34533
rect 9309 34524 9321 34527
rect 8904 34496 9321 34524
rect 8904 34484 8910 34496
rect 9309 34493 9321 34496
rect 9355 34493 9367 34527
rect 9309 34487 9367 34493
rect 16485 34527 16543 34533
rect 16485 34493 16497 34527
rect 16531 34524 16543 34527
rect 17770 34524 17776 34536
rect 16531 34496 17776 34524
rect 16531 34493 16543 34496
rect 16485 34487 16543 34493
rect 17770 34484 17776 34496
rect 17828 34484 17834 34536
rect 18892 34524 18920 34552
rect 18892 34496 19564 34524
rect 19061 34459 19119 34465
rect 19061 34425 19073 34459
rect 19107 34456 19119 34459
rect 19334 34456 19340 34468
rect 19107 34428 19340 34456
rect 19107 34425 19119 34428
rect 19061 34419 19119 34425
rect 19334 34416 19340 34428
rect 19392 34416 19398 34468
rect 19536 34456 19564 34496
rect 19610 34484 19616 34536
rect 19668 34484 19674 34536
rect 20165 34527 20223 34533
rect 20165 34493 20177 34527
rect 20211 34493 20223 34527
rect 20901 34527 20959 34533
rect 20901 34524 20913 34527
rect 20165 34487 20223 34493
rect 20272 34496 20913 34524
rect 20180 34456 20208 34487
rect 19536 34428 20208 34456
rect 15010 34348 15016 34400
rect 15068 34388 15074 34400
rect 15105 34391 15163 34397
rect 15105 34388 15117 34391
rect 15068 34360 15117 34388
rect 15068 34348 15074 34360
rect 15105 34357 15117 34360
rect 15151 34357 15163 34391
rect 15105 34351 15163 34357
rect 19518 34348 19524 34400
rect 19576 34388 19582 34400
rect 20272 34388 20300 34496
rect 20901 34493 20913 34496
rect 20947 34524 20959 34527
rect 21284 34524 21312 34555
rect 20947 34496 21312 34524
rect 21468 34524 21496 34555
rect 22002 34552 22008 34604
rect 22060 34552 22066 34604
rect 22296 34601 22324 34632
rect 22922 34620 22928 34672
rect 22980 34660 22986 34672
rect 23753 34663 23811 34669
rect 23753 34660 23765 34663
rect 22980 34632 23765 34660
rect 22980 34620 22986 34632
rect 23753 34629 23765 34632
rect 23799 34629 23811 34663
rect 23753 34623 23811 34629
rect 23845 34663 23903 34669
rect 23845 34629 23857 34663
rect 23891 34660 23903 34663
rect 24302 34660 24308 34672
rect 23891 34632 24308 34660
rect 23891 34629 23903 34632
rect 23845 34623 23903 34629
rect 24302 34620 24308 34632
rect 24360 34660 24366 34672
rect 24765 34663 24823 34669
rect 24765 34660 24777 34663
rect 24360 34632 24777 34660
rect 24360 34620 24366 34632
rect 24765 34629 24777 34632
rect 24811 34629 24823 34663
rect 24765 34623 24823 34629
rect 26786 34620 26792 34672
rect 26844 34620 26850 34672
rect 27709 34663 27767 34669
rect 27709 34660 27721 34663
rect 26896 34632 27721 34660
rect 22189 34595 22247 34601
rect 22189 34592 22201 34595
rect 22112 34564 22201 34592
rect 22112 34536 22140 34564
rect 22189 34561 22201 34564
rect 22235 34561 22247 34595
rect 22189 34555 22247 34561
rect 22281 34595 22339 34601
rect 22281 34561 22293 34595
rect 22327 34561 22339 34595
rect 22281 34555 22339 34561
rect 22557 34595 22615 34601
rect 22557 34561 22569 34595
rect 22603 34561 22615 34595
rect 22557 34555 22615 34561
rect 22741 34595 22799 34601
rect 22741 34561 22753 34595
rect 22787 34592 22799 34595
rect 23477 34595 23535 34601
rect 23477 34592 23489 34595
rect 22787 34564 23489 34592
rect 22787 34561 22799 34564
rect 22741 34555 22799 34561
rect 23477 34561 23489 34564
rect 23523 34561 23535 34595
rect 23477 34555 23535 34561
rect 23570 34595 23628 34601
rect 23570 34561 23582 34595
rect 23616 34592 23628 34595
rect 23658 34592 23664 34604
rect 23616 34564 23664 34592
rect 23616 34561 23628 34564
rect 23570 34555 23628 34561
rect 22094 34524 22100 34536
rect 21468 34496 22100 34524
rect 20947 34493 20959 34496
rect 20901 34487 20959 34493
rect 22094 34484 22100 34496
rect 22152 34484 22158 34536
rect 22373 34527 22431 34533
rect 22373 34493 22385 34527
rect 22419 34493 22431 34527
rect 22572 34524 22600 34555
rect 23584 34524 23612 34555
rect 23658 34552 23664 34564
rect 23716 34552 23722 34604
rect 23983 34595 24041 34601
rect 23983 34561 23995 34595
rect 24029 34592 24041 34595
rect 24581 34595 24639 34601
rect 24581 34592 24593 34595
rect 24029 34564 24593 34592
rect 24029 34561 24041 34564
rect 23983 34555 24041 34561
rect 24581 34561 24593 34564
rect 24627 34561 24639 34595
rect 24581 34555 24639 34561
rect 26329 34595 26387 34601
rect 26329 34561 26341 34595
rect 26375 34592 26387 34595
rect 26510 34592 26516 34604
rect 26375 34564 26516 34592
rect 26375 34561 26387 34564
rect 26329 34555 26387 34561
rect 22572 34496 23612 34524
rect 24596 34524 24624 34555
rect 26510 34552 26516 34564
rect 26568 34552 26574 34604
rect 26697 34595 26755 34601
rect 26697 34561 26709 34595
rect 26743 34592 26755 34595
rect 26896 34592 26924 34632
rect 27709 34629 27721 34632
rect 27755 34629 27767 34663
rect 27709 34623 27767 34629
rect 26743 34564 26924 34592
rect 26743 34561 26755 34564
rect 26697 34555 26755 34561
rect 26970 34552 26976 34604
rect 27028 34552 27034 34604
rect 27157 34595 27215 34601
rect 27157 34561 27169 34595
rect 27203 34561 27215 34595
rect 27157 34555 27215 34561
rect 24854 34524 24860 34536
rect 24596 34496 24860 34524
rect 22373 34487 22431 34493
rect 22388 34456 22416 34487
rect 24854 34484 24860 34496
rect 24912 34484 24918 34536
rect 25590 34484 25596 34536
rect 25648 34524 25654 34536
rect 27172 34524 27200 34555
rect 27430 34552 27436 34604
rect 27488 34592 27494 34604
rect 27525 34595 27583 34601
rect 27525 34592 27537 34595
rect 27488 34564 27537 34592
rect 27488 34552 27494 34564
rect 27525 34561 27537 34564
rect 27571 34561 27583 34595
rect 27525 34555 27583 34561
rect 25648 34496 27200 34524
rect 25648 34484 25654 34496
rect 27246 34484 27252 34536
rect 27304 34484 27310 34536
rect 27341 34527 27399 34533
rect 27341 34493 27353 34527
rect 27387 34524 27399 34527
rect 27982 34524 27988 34536
rect 27387 34496 27988 34524
rect 27387 34493 27399 34496
rect 27341 34487 27399 34493
rect 27982 34484 27988 34496
rect 28040 34484 28046 34536
rect 22922 34456 22928 34468
rect 22388 34428 22928 34456
rect 22922 34416 22928 34428
rect 22980 34416 22986 34468
rect 26602 34416 26608 34468
rect 26660 34416 26666 34468
rect 19576 34360 20300 34388
rect 24949 34391 25007 34397
rect 19576 34348 19582 34360
rect 24949 34357 24961 34391
rect 24995 34388 25007 34391
rect 25406 34388 25412 34400
rect 24995 34360 25412 34388
rect 24995 34357 25007 34360
rect 24949 34351 25007 34357
rect 25406 34348 25412 34360
rect 25464 34348 25470 34400
rect 1104 34298 28888 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 28888 34298
rect 1104 34224 28888 34246
rect 16206 34144 16212 34196
rect 16264 34144 16270 34196
rect 17770 34144 17776 34196
rect 17828 34184 17834 34196
rect 23109 34187 23167 34193
rect 17828 34156 20668 34184
rect 17828 34144 17834 34156
rect 18049 34119 18107 34125
rect 18049 34085 18061 34119
rect 18095 34116 18107 34119
rect 18690 34116 18696 34128
rect 18095 34088 18696 34116
rect 18095 34085 18107 34088
rect 18049 34079 18107 34085
rect 18690 34076 18696 34088
rect 18748 34076 18754 34128
rect 17494 34048 17500 34060
rect 15764 34020 17500 34048
rect 15010 33940 15016 33992
rect 15068 33980 15074 33992
rect 15764 33989 15792 34020
rect 17494 34008 17500 34020
rect 17552 34008 17558 34060
rect 18417 34051 18475 34057
rect 18417 34048 18429 34051
rect 17972 34020 18429 34048
rect 15749 33983 15807 33989
rect 15749 33980 15761 33983
rect 15068 33952 15761 33980
rect 15068 33940 15074 33952
rect 15749 33949 15761 33952
rect 15795 33949 15807 33983
rect 15749 33943 15807 33949
rect 16025 33983 16083 33989
rect 16025 33949 16037 33983
rect 16071 33949 16083 33983
rect 16025 33943 16083 33949
rect 16209 33983 16267 33989
rect 16209 33949 16221 33983
rect 16255 33980 16267 33983
rect 16666 33980 16672 33992
rect 16255 33952 16672 33980
rect 16255 33949 16267 33952
rect 16209 33943 16267 33949
rect 15102 33872 15108 33924
rect 15160 33912 15166 33924
rect 15565 33915 15623 33921
rect 15565 33912 15577 33915
rect 15160 33884 15577 33912
rect 15160 33872 15166 33884
rect 15565 33881 15577 33884
rect 15611 33881 15623 33915
rect 16040 33912 16068 33943
rect 16666 33940 16672 33952
rect 16724 33940 16730 33992
rect 17972 33989 18000 34020
rect 18417 34017 18429 34020
rect 18463 34017 18475 34051
rect 18417 34011 18475 34017
rect 18598 34008 18604 34060
rect 18656 34048 18662 34060
rect 18969 34051 19027 34057
rect 18969 34048 18981 34051
rect 18656 34020 18981 34048
rect 18656 34008 18662 34020
rect 18969 34017 18981 34020
rect 19015 34048 19027 34051
rect 19150 34048 19156 34060
rect 19015 34020 19156 34048
rect 19015 34017 19027 34020
rect 18969 34011 19027 34017
rect 19150 34008 19156 34020
rect 19208 34008 19214 34060
rect 20640 34057 20668 34156
rect 23109 34153 23121 34187
rect 23155 34184 23167 34187
rect 23198 34184 23204 34196
rect 23155 34156 23204 34184
rect 23155 34153 23167 34156
rect 23109 34147 23167 34153
rect 20625 34051 20683 34057
rect 20625 34017 20637 34051
rect 20671 34017 20683 34051
rect 20625 34011 20683 34017
rect 21729 34051 21787 34057
rect 21729 34017 21741 34051
rect 21775 34048 21787 34051
rect 22094 34048 22100 34060
rect 21775 34020 22100 34048
rect 21775 34017 21787 34020
rect 21729 34011 21787 34017
rect 17773 33983 17831 33989
rect 17773 33949 17785 33983
rect 17819 33949 17831 33983
rect 17773 33943 17831 33949
rect 17957 33983 18015 33989
rect 17957 33949 17969 33983
rect 18003 33949 18015 33983
rect 18325 33983 18383 33989
rect 18325 33980 18337 33983
rect 17957 33943 18015 33949
rect 18156 33952 18337 33980
rect 17788 33912 17816 33943
rect 18046 33912 18052 33924
rect 16040 33884 18052 33912
rect 15565 33875 15623 33881
rect 18046 33872 18052 33884
rect 18104 33872 18110 33924
rect 15930 33804 15936 33856
rect 15988 33804 15994 33856
rect 17862 33804 17868 33856
rect 17920 33804 17926 33856
rect 18156 33844 18184 33952
rect 18325 33949 18337 33952
rect 18371 33949 18383 33983
rect 18325 33943 18383 33949
rect 18233 33915 18291 33921
rect 18233 33881 18245 33915
rect 18279 33912 18291 33915
rect 18616 33912 18644 34008
rect 20640 33980 20668 34011
rect 22094 34008 22100 34020
rect 22152 34048 22158 34060
rect 22833 34051 22891 34057
rect 22833 34048 22845 34051
rect 22152 34020 22845 34048
rect 22152 34008 22158 34020
rect 22833 34017 22845 34020
rect 22879 34048 22891 34051
rect 23124 34048 23152 34147
rect 23198 34144 23204 34156
rect 23256 34144 23262 34196
rect 25777 34187 25835 34193
rect 25777 34153 25789 34187
rect 25823 34184 25835 34187
rect 26970 34184 26976 34196
rect 25823 34156 26976 34184
rect 25823 34153 25835 34156
rect 25777 34147 25835 34153
rect 26970 34144 26976 34156
rect 27028 34144 27034 34196
rect 22879 34020 23152 34048
rect 22879 34017 22891 34020
rect 22833 34011 22891 34017
rect 27982 34008 27988 34060
rect 28040 34008 28046 34060
rect 20717 33983 20775 33989
rect 20717 33980 20729 33983
rect 20640 33952 20729 33980
rect 20717 33949 20729 33952
rect 20763 33980 20775 33983
rect 21174 33980 21180 33992
rect 20763 33952 21180 33980
rect 20763 33949 20775 33952
rect 20717 33943 20775 33949
rect 21174 33940 21180 33952
rect 21232 33940 21238 33992
rect 21266 33940 21272 33992
rect 21324 33980 21330 33992
rect 21913 33983 21971 33989
rect 21913 33980 21925 33983
rect 21324 33952 21925 33980
rect 21324 33940 21330 33952
rect 21913 33949 21925 33952
rect 21959 33980 21971 33983
rect 21959 33952 22600 33980
rect 21959 33949 21971 33952
rect 21913 33943 21971 33949
rect 18279 33884 18644 33912
rect 18279 33881 18291 33884
rect 18233 33875 18291 33881
rect 19978 33872 19984 33924
rect 20036 33912 20042 33924
rect 20358 33915 20416 33921
rect 20358 33912 20370 33915
rect 20036 33884 20370 33912
rect 20036 33872 20042 33884
rect 20358 33881 20370 33884
rect 20404 33881 20416 33915
rect 20358 33875 20416 33881
rect 22097 33915 22155 33921
rect 22097 33881 22109 33915
rect 22143 33912 22155 33915
rect 22462 33912 22468 33924
rect 22143 33884 22468 33912
rect 22143 33881 22155 33884
rect 22097 33875 22155 33881
rect 22462 33872 22468 33884
rect 22520 33872 22526 33924
rect 18874 33844 18880 33856
rect 18156 33816 18880 33844
rect 18874 33804 18880 33816
rect 18932 33844 18938 33856
rect 19242 33844 19248 33856
rect 18932 33816 19248 33844
rect 18932 33804 18938 33816
rect 19242 33804 19248 33816
rect 19300 33804 19306 33856
rect 22189 33847 22247 33853
rect 22189 33813 22201 33847
rect 22235 33844 22247 33847
rect 22278 33844 22284 33856
rect 22235 33816 22284 33844
rect 22235 33813 22247 33816
rect 22189 33807 22247 33813
rect 22278 33804 22284 33816
rect 22336 33804 22342 33856
rect 22572 33844 22600 33952
rect 25222 33940 25228 33992
rect 25280 33940 25286 33992
rect 25406 33940 25412 33992
rect 25464 33940 25470 33992
rect 25590 33940 25596 33992
rect 25648 33940 25654 33992
rect 22922 33872 22928 33924
rect 22980 33872 22986 33924
rect 25501 33915 25559 33921
rect 25501 33881 25513 33915
rect 25547 33912 25559 33915
rect 27246 33912 27252 33924
rect 25547 33884 27252 33912
rect 25547 33881 25559 33884
rect 25501 33875 25559 33881
rect 27246 33872 27252 33884
rect 27304 33872 27310 33924
rect 23125 33847 23183 33853
rect 23125 33844 23137 33847
rect 22572 33816 23137 33844
rect 23125 33813 23137 33816
rect 23171 33813 23183 33847
rect 23125 33807 23183 33813
rect 23293 33847 23351 33853
rect 23293 33813 23305 33847
rect 23339 33844 23351 33847
rect 24026 33844 24032 33856
rect 23339 33816 24032 33844
rect 23339 33813 23351 33816
rect 23293 33807 23351 33813
rect 24026 33804 24032 33816
rect 24084 33804 24090 33856
rect 26510 33804 26516 33856
rect 26568 33844 26574 33856
rect 27433 33847 27491 33853
rect 27433 33844 27445 33847
rect 26568 33816 27445 33844
rect 26568 33804 26574 33816
rect 27433 33813 27445 33816
rect 27479 33813 27491 33847
rect 27433 33807 27491 33813
rect 1104 33754 28888 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 28888 33754
rect 1104 33680 28888 33702
rect 3697 33643 3755 33649
rect 3697 33609 3709 33643
rect 3743 33640 3755 33643
rect 4614 33640 4620 33652
rect 3743 33612 4620 33640
rect 3743 33609 3755 33612
rect 3697 33603 3755 33609
rect 4614 33600 4620 33612
rect 4672 33600 4678 33652
rect 15933 33643 15991 33649
rect 15933 33609 15945 33643
rect 15979 33609 15991 33643
rect 15933 33603 15991 33609
rect 15289 33575 15347 33581
rect 15289 33541 15301 33575
rect 15335 33572 15347 33575
rect 15470 33572 15476 33584
rect 15335 33544 15476 33572
rect 15335 33541 15347 33544
rect 15289 33535 15347 33541
rect 15470 33532 15476 33544
rect 15528 33572 15534 33584
rect 15948 33572 15976 33603
rect 16666 33600 16672 33652
rect 16724 33600 16730 33652
rect 17037 33643 17095 33649
rect 17037 33609 17049 33643
rect 17083 33640 17095 33643
rect 17586 33640 17592 33652
rect 17083 33612 17592 33640
rect 17083 33609 17095 33612
rect 17037 33603 17095 33609
rect 17586 33600 17592 33612
rect 17644 33600 17650 33652
rect 19150 33600 19156 33652
rect 19208 33640 19214 33652
rect 19208 33612 19472 33640
rect 19208 33600 19214 33612
rect 17129 33575 17187 33581
rect 17129 33572 17141 33575
rect 15528 33544 15792 33572
rect 15948 33544 17141 33572
rect 15528 33532 15534 33544
rect 3510 33464 3516 33516
rect 3568 33464 3574 33516
rect 12796 33507 12854 33513
rect 12796 33473 12808 33507
rect 12842 33504 12854 33507
rect 13262 33504 13268 33516
rect 12842 33476 13268 33504
rect 12842 33473 12854 33476
rect 12796 33467 12854 33473
rect 13262 33464 13268 33476
rect 13320 33464 13326 33516
rect 15010 33464 15016 33516
rect 15068 33464 15074 33516
rect 15102 33464 15108 33516
rect 15160 33504 15166 33516
rect 15565 33507 15623 33513
rect 15160 33476 15205 33504
rect 15160 33464 15166 33476
rect 15565 33473 15577 33507
rect 15611 33473 15623 33507
rect 15764 33504 15792 33544
rect 17129 33541 17141 33544
rect 17175 33541 17187 33575
rect 17129 33535 17187 33541
rect 17862 33532 17868 33584
rect 17920 33572 17926 33584
rect 18018 33575 18076 33581
rect 18018 33572 18030 33575
rect 17920 33544 18030 33572
rect 17920 33532 17926 33544
rect 18018 33541 18030 33544
rect 18064 33541 18076 33575
rect 18018 33535 18076 33541
rect 18138 33532 18144 33584
rect 18196 33572 18202 33584
rect 19444 33581 19472 33612
rect 21174 33600 21180 33652
rect 21232 33600 21238 33652
rect 23198 33600 23204 33652
rect 23256 33600 23262 33652
rect 19429 33575 19487 33581
rect 18196 33544 18828 33572
rect 18196 33532 18202 33544
rect 16485 33507 16543 33513
rect 16485 33504 16497 33507
rect 15764 33476 16497 33504
rect 15565 33467 15623 33473
rect 16485 33473 16497 33476
rect 16531 33473 16543 33507
rect 16485 33467 16543 33473
rect 2958 33396 2964 33448
rect 3016 33436 3022 33448
rect 3329 33439 3387 33445
rect 3329 33436 3341 33439
rect 3016 33408 3341 33436
rect 3016 33396 3022 33408
rect 3329 33405 3341 33408
rect 3375 33405 3387 33439
rect 3329 33399 3387 33405
rect 8846 33396 8852 33448
rect 8904 33436 8910 33448
rect 12529 33439 12587 33445
rect 12529 33436 12541 33439
rect 8904 33408 12541 33436
rect 8904 33396 8910 33408
rect 12529 33405 12541 33408
rect 12575 33405 12587 33439
rect 12529 33399 12587 33405
rect 14553 33439 14611 33445
rect 14553 33405 14565 33439
rect 14599 33405 14611 33439
rect 14553 33399 14611 33405
rect 13906 33328 13912 33380
rect 13964 33368 13970 33380
rect 14568 33368 14596 33399
rect 15286 33396 15292 33448
rect 15344 33436 15350 33448
rect 15473 33439 15531 33445
rect 15473 33436 15485 33439
rect 15344 33408 15485 33436
rect 15344 33396 15350 33408
rect 15473 33405 15485 33408
rect 15519 33405 15531 33439
rect 15580 33436 15608 33467
rect 17494 33464 17500 33516
rect 17552 33464 17558 33516
rect 17770 33464 17776 33516
rect 17828 33464 17834 33516
rect 16025 33439 16083 33445
rect 16025 33436 16037 33439
rect 15580 33408 16037 33436
rect 15473 33399 15531 33405
rect 16025 33405 16037 33408
rect 16071 33405 16083 33439
rect 16025 33399 16083 33405
rect 17218 33396 17224 33448
rect 17276 33396 17282 33448
rect 18800 33436 18828 33544
rect 19429 33541 19441 33575
rect 19475 33541 19487 33575
rect 19629 33575 19687 33581
rect 19629 33572 19641 33575
rect 19429 33535 19487 33541
rect 19536 33544 19641 33572
rect 19242 33464 19248 33516
rect 19300 33504 19306 33516
rect 19536 33504 19564 33544
rect 19629 33541 19641 33544
rect 19675 33541 19687 33575
rect 19629 33535 19687 33541
rect 19886 33532 19892 33584
rect 19944 33532 19950 33584
rect 22094 33513 22100 33516
rect 19300 33476 19564 33504
rect 19300 33464 19306 33476
rect 22088 33467 22100 33513
rect 22094 33464 22100 33467
rect 22152 33464 22158 33516
rect 22462 33464 22468 33516
rect 22520 33504 22526 33516
rect 23293 33507 23351 33513
rect 23293 33504 23305 33507
rect 22520 33476 23305 33504
rect 22520 33464 22526 33476
rect 23293 33473 23305 33476
rect 23339 33473 23351 33507
rect 23293 33467 23351 33473
rect 23477 33507 23535 33513
rect 23477 33473 23489 33507
rect 23523 33504 23535 33507
rect 26602 33504 26608 33516
rect 23523 33476 26608 33504
rect 23523 33473 23535 33476
rect 23477 33467 23535 33473
rect 26602 33464 26608 33476
rect 26660 33464 26666 33516
rect 20990 33436 20996 33448
rect 18800 33408 20996 33436
rect 20990 33396 20996 33408
rect 21048 33396 21054 33448
rect 21174 33396 21180 33448
rect 21232 33436 21238 33448
rect 21821 33439 21879 33445
rect 21821 33436 21833 33439
rect 21232 33408 21833 33436
rect 21232 33396 21238 33408
rect 21821 33405 21833 33408
rect 21867 33405 21879 33439
rect 21821 33399 21879 33405
rect 13964 33340 14596 33368
rect 13964 33328 13970 33340
rect 15378 33328 15384 33380
rect 15436 33368 15442 33380
rect 15930 33368 15936 33380
rect 15436 33340 15936 33368
rect 15436 33328 15442 33340
rect 15930 33328 15936 33340
rect 15988 33368 15994 33380
rect 16117 33371 16175 33377
rect 16117 33368 16129 33371
rect 15988 33340 16129 33368
rect 15988 33328 15994 33340
rect 16117 33337 16129 33340
rect 16163 33337 16175 33371
rect 16117 33331 16175 33337
rect 13998 33260 14004 33312
rect 14056 33260 14062 33312
rect 19518 33260 19524 33312
rect 19576 33300 19582 33312
rect 19613 33303 19671 33309
rect 19613 33300 19625 33303
rect 19576 33272 19625 33300
rect 19576 33260 19582 33272
rect 19613 33269 19625 33272
rect 19659 33269 19671 33303
rect 19613 33263 19671 33269
rect 19797 33303 19855 33309
rect 19797 33269 19809 33303
rect 19843 33300 19855 33303
rect 21266 33300 21272 33312
rect 19843 33272 21272 33300
rect 19843 33269 19855 33272
rect 19797 33263 19855 33269
rect 21266 33260 21272 33272
rect 21324 33260 21330 33312
rect 23290 33260 23296 33312
rect 23348 33260 23354 33312
rect 1104 33210 28888 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 28888 33210
rect 1104 33136 28888 33158
rect 1581 33099 1639 33105
rect 1581 33065 1593 33099
rect 1627 33096 1639 33099
rect 3510 33096 3516 33108
rect 1627 33068 3516 33096
rect 1627 33065 1639 33068
rect 1581 33059 1639 33065
rect 3510 33056 3516 33068
rect 3568 33056 3574 33108
rect 13262 33056 13268 33108
rect 13320 33056 13326 33108
rect 13541 33099 13599 33105
rect 13541 33065 13553 33099
rect 13587 33065 13599 33099
rect 13541 33059 13599 33065
rect 12526 32988 12532 33040
rect 12584 33028 12590 33040
rect 13556 33028 13584 33059
rect 13630 33056 13636 33108
rect 13688 33096 13694 33108
rect 15102 33096 15108 33108
rect 13688 33068 15108 33096
rect 13688 33056 13694 33068
rect 15102 33056 15108 33068
rect 15160 33056 15166 33108
rect 18509 33099 18567 33105
rect 18509 33065 18521 33099
rect 18555 33096 18567 33099
rect 19610 33096 19616 33108
rect 18555 33068 19616 33096
rect 18555 33065 18567 33068
rect 18509 33059 18567 33065
rect 19610 33056 19616 33068
rect 19668 33056 19674 33108
rect 21266 33056 21272 33108
rect 21324 33056 21330 33108
rect 21637 33099 21695 33105
rect 21637 33065 21649 33099
rect 21683 33096 21695 33099
rect 22094 33096 22100 33108
rect 21683 33068 22100 33096
rect 21683 33065 21695 33068
rect 21637 33059 21695 33065
rect 22094 33056 22100 33068
rect 22152 33056 22158 33108
rect 22922 33056 22928 33108
rect 22980 33096 22986 33108
rect 23201 33099 23259 33105
rect 23201 33096 23213 33099
rect 22980 33068 23213 33096
rect 22980 33056 22986 33068
rect 23201 33065 23213 33068
rect 23247 33065 23259 33099
rect 23201 33059 23259 33065
rect 14090 33028 14096 33040
rect 12584 33000 14096 33028
rect 12584 32988 12590 33000
rect 14090 32988 14096 33000
rect 14148 32988 14154 33040
rect 21174 32988 21180 33040
rect 21232 32988 21238 33040
rect 12345 32963 12403 32969
rect 12345 32929 12357 32963
rect 12391 32960 12403 32963
rect 12805 32963 12863 32969
rect 12805 32960 12817 32963
rect 12391 32932 12817 32960
rect 12391 32929 12403 32932
rect 12345 32923 12403 32929
rect 12805 32929 12817 32932
rect 12851 32929 12863 32963
rect 12805 32923 12863 32929
rect 12894 32920 12900 32972
rect 12952 32960 12958 32972
rect 16574 32960 16580 32972
rect 12952 32932 16580 32960
rect 12952 32920 12958 32932
rect 16574 32920 16580 32932
rect 16632 32960 16638 32972
rect 17218 32960 17224 32972
rect 16632 32932 17224 32960
rect 16632 32920 16638 32932
rect 17218 32920 17224 32932
rect 17276 32920 17282 32972
rect 18417 32963 18475 32969
rect 18417 32929 18429 32963
rect 18463 32960 18475 32963
rect 18598 32960 18604 32972
rect 18463 32932 18604 32960
rect 18463 32929 18475 32932
rect 18417 32923 18475 32929
rect 18598 32920 18604 32932
rect 18656 32920 18662 32972
rect 20993 32963 21051 32969
rect 20993 32929 21005 32963
rect 21039 32960 21051 32963
rect 21192 32960 21220 32988
rect 21818 32960 21824 32972
rect 21039 32932 21824 32960
rect 21039 32929 21051 32932
rect 20993 32923 21051 32929
rect 21818 32920 21824 32932
rect 21876 32920 21882 32972
rect 23216 32960 23244 33059
rect 24854 33056 24860 33108
rect 24912 33096 24918 33108
rect 25225 33099 25283 33105
rect 25225 33096 25237 33099
rect 24912 33068 25237 33096
rect 24912 33056 24918 33068
rect 25225 33065 25237 33068
rect 25271 33065 25283 33099
rect 25225 33059 25283 33065
rect 25409 33031 25467 33037
rect 25409 32997 25421 33031
rect 25455 32997 25467 33031
rect 25409 32991 25467 32997
rect 23845 32963 23903 32969
rect 23845 32960 23857 32963
rect 23216 32932 23857 32960
rect 23845 32929 23857 32932
rect 23891 32929 23903 32963
rect 23845 32923 23903 32929
rect 24044 32932 24716 32960
rect 24044 32904 24072 32932
rect 842 32852 848 32904
rect 900 32892 906 32904
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 900 32864 1409 32892
rect 900 32852 906 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 11882 32852 11888 32904
rect 11940 32892 11946 32904
rect 12253 32895 12311 32901
rect 12253 32892 12265 32895
rect 11940 32864 12265 32892
rect 11940 32852 11946 32864
rect 12253 32861 12265 32864
rect 12299 32861 12311 32895
rect 12253 32855 12311 32861
rect 12434 32852 12440 32904
rect 12492 32852 12498 32904
rect 12529 32895 12587 32901
rect 12529 32861 12541 32895
rect 12575 32892 12587 32895
rect 12618 32892 12624 32904
rect 12575 32864 12624 32892
rect 12575 32861 12587 32864
rect 12529 32855 12587 32861
rect 12618 32852 12624 32864
rect 12676 32852 12682 32904
rect 12713 32895 12771 32901
rect 12713 32861 12725 32895
rect 12759 32861 12771 32895
rect 12713 32855 12771 32861
rect 13081 32895 13139 32901
rect 13081 32861 13093 32895
rect 13127 32892 13139 32895
rect 13998 32892 14004 32904
rect 13127 32864 14004 32892
rect 13127 32861 13139 32864
rect 13081 32855 13139 32861
rect 12728 32824 12756 32855
rect 13998 32852 14004 32864
rect 14056 32852 14062 32904
rect 15286 32852 15292 32904
rect 15344 32852 15350 32904
rect 15378 32852 15384 32904
rect 15436 32852 15442 32904
rect 15470 32852 15476 32904
rect 15528 32892 15534 32904
rect 15565 32895 15623 32901
rect 15565 32892 15577 32895
rect 15528 32864 15577 32892
rect 15528 32852 15534 32864
rect 15565 32861 15577 32864
rect 15611 32861 15623 32895
rect 15565 32855 15623 32861
rect 18690 32852 18696 32904
rect 18748 32852 18754 32904
rect 21177 32895 21235 32901
rect 21177 32861 21189 32895
rect 21223 32861 21235 32895
rect 21177 32855 21235 32861
rect 21453 32895 21511 32901
rect 21453 32861 21465 32895
rect 21499 32892 21511 32895
rect 23290 32892 23296 32904
rect 21499 32864 23296 32892
rect 21499 32861 21511 32864
rect 21453 32855 21511 32861
rect 13725 32827 13783 32833
rect 12728 32796 13400 32824
rect 13372 32765 13400 32796
rect 13725 32793 13737 32827
rect 13771 32824 13783 32827
rect 14182 32824 14188 32836
rect 13771 32796 14188 32824
rect 13771 32793 13783 32796
rect 13725 32787 13783 32793
rect 14182 32784 14188 32796
rect 14240 32784 14246 32836
rect 20714 32784 20720 32836
rect 20772 32833 20778 32836
rect 20772 32824 20784 32833
rect 20772 32796 20817 32824
rect 20772 32787 20784 32796
rect 20772 32784 20778 32787
rect 13357 32759 13415 32765
rect 13357 32725 13369 32759
rect 13403 32725 13415 32759
rect 13357 32719 13415 32725
rect 13525 32759 13583 32765
rect 13525 32725 13537 32759
rect 13571 32756 13583 32759
rect 13814 32756 13820 32768
rect 13571 32728 13820 32756
rect 13571 32725 13583 32728
rect 13525 32719 13583 32725
rect 13814 32716 13820 32728
rect 13872 32716 13878 32768
rect 15562 32716 15568 32768
rect 15620 32756 15626 32768
rect 15749 32759 15807 32765
rect 15749 32756 15761 32759
rect 15620 32728 15761 32756
rect 15620 32716 15626 32728
rect 15749 32725 15761 32728
rect 15795 32725 15807 32759
rect 15749 32719 15807 32725
rect 18877 32759 18935 32765
rect 18877 32725 18889 32759
rect 18923 32756 18935 32759
rect 19242 32756 19248 32768
rect 18923 32728 19248 32756
rect 18923 32725 18935 32728
rect 18877 32719 18935 32725
rect 19242 32716 19248 32728
rect 19300 32716 19306 32768
rect 19518 32716 19524 32768
rect 19576 32756 19582 32768
rect 19613 32759 19671 32765
rect 19613 32756 19625 32759
rect 19576 32728 19625 32756
rect 19576 32716 19582 32728
rect 19613 32725 19625 32728
rect 19659 32725 19671 32759
rect 21192 32756 21220 32855
rect 23290 32852 23296 32864
rect 23348 32852 23354 32904
rect 24026 32852 24032 32904
rect 24084 32852 24090 32904
rect 24213 32895 24271 32901
rect 24213 32861 24225 32895
rect 24259 32892 24271 32895
rect 24302 32892 24308 32904
rect 24259 32864 24308 32892
rect 24259 32861 24271 32864
rect 24213 32855 24271 32861
rect 24302 32852 24308 32864
rect 24360 32852 24366 32904
rect 24688 32901 24716 32932
rect 24854 32920 24860 32972
rect 24912 32920 24918 32972
rect 24673 32895 24731 32901
rect 24673 32861 24685 32895
rect 24719 32861 24731 32895
rect 25424 32892 25452 32991
rect 27617 32963 27675 32969
rect 27617 32960 27629 32963
rect 26712 32932 27629 32960
rect 26142 32892 26148 32904
rect 25424 32864 26148 32892
rect 24673 32855 24731 32861
rect 22088 32827 22146 32833
rect 22088 32793 22100 32827
rect 22134 32824 22146 32827
rect 22186 32824 22192 32836
rect 22134 32796 22192 32824
rect 22134 32793 22146 32796
rect 22088 32787 22146 32793
rect 22186 32784 22192 32796
rect 22244 32784 22250 32836
rect 22370 32784 22376 32836
rect 22428 32824 22434 32836
rect 24121 32827 24179 32833
rect 24121 32824 24133 32827
rect 22428 32796 24133 32824
rect 22428 32784 22434 32796
rect 24121 32793 24133 32796
rect 24167 32793 24179 32827
rect 24121 32787 24179 32793
rect 22278 32756 22284 32768
rect 21192 32728 22284 32756
rect 19613 32719 19671 32725
rect 22278 32716 22284 32728
rect 22336 32716 22342 32768
rect 23290 32716 23296 32768
rect 23348 32716 23354 32768
rect 24210 32716 24216 32768
rect 24268 32756 24274 32768
rect 24489 32759 24547 32765
rect 24489 32756 24501 32759
rect 24268 32728 24501 32756
rect 24268 32716 24274 32728
rect 24489 32725 24501 32728
rect 24535 32725 24547 32759
rect 24688 32756 24716 32855
rect 26142 32852 26148 32864
rect 26200 32892 26206 32904
rect 26712 32901 26740 32932
rect 27617 32929 27629 32932
rect 27663 32929 27675 32963
rect 27617 32923 27675 32929
rect 27982 32920 27988 32972
rect 28040 32960 28046 32972
rect 28169 32963 28227 32969
rect 28169 32960 28181 32963
rect 28040 32932 28181 32960
rect 28040 32920 28046 32932
rect 28169 32929 28181 32932
rect 28215 32929 28227 32963
rect 28169 32923 28227 32929
rect 26605 32895 26663 32901
rect 26605 32892 26617 32895
rect 26200 32864 26617 32892
rect 26200 32852 26206 32864
rect 26605 32861 26617 32864
rect 26651 32861 26663 32895
rect 26605 32855 26663 32861
rect 26697 32895 26755 32901
rect 26697 32861 26709 32895
rect 26743 32861 26755 32895
rect 26697 32855 26755 32861
rect 26786 32852 26792 32904
rect 26844 32892 26850 32904
rect 26973 32895 27031 32901
rect 26973 32892 26985 32895
rect 26844 32864 26985 32892
rect 26844 32852 26850 32864
rect 26973 32861 26985 32864
rect 27019 32861 27031 32895
rect 26973 32855 27031 32861
rect 25041 32827 25099 32833
rect 25041 32793 25053 32827
rect 25087 32824 25099 32827
rect 25590 32824 25596 32836
rect 25087 32796 25596 32824
rect 25087 32793 25099 32796
rect 25041 32787 25099 32793
rect 25590 32784 25596 32796
rect 25648 32784 25654 32836
rect 25682 32784 25688 32836
rect 25740 32824 25746 32836
rect 26881 32827 26939 32833
rect 26881 32824 26893 32827
rect 25740 32796 26893 32824
rect 25740 32784 25746 32796
rect 26881 32793 26893 32796
rect 26927 32793 26939 32827
rect 26881 32787 26939 32793
rect 24762 32756 24768 32768
rect 24688 32728 24768 32756
rect 24489 32719 24547 32725
rect 24762 32716 24768 32728
rect 24820 32756 24826 32768
rect 26786 32765 26792 32768
rect 25241 32759 25299 32765
rect 25241 32756 25253 32759
rect 24820 32728 25253 32756
rect 24820 32716 24826 32728
rect 25241 32725 25253 32728
rect 25287 32725 25299 32759
rect 25241 32719 25299 32725
rect 26782 32719 26792 32765
rect 26786 32716 26792 32719
rect 26844 32716 26850 32768
rect 26896 32756 26924 32787
rect 27157 32759 27215 32765
rect 27157 32756 27169 32759
rect 26896 32728 27169 32756
rect 27157 32725 27169 32728
rect 27203 32725 27215 32759
rect 27157 32719 27215 32725
rect 1104 32666 28888 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 28888 32666
rect 1104 32592 28888 32614
rect 12621 32555 12679 32561
rect 12621 32521 12633 32555
rect 12667 32552 12679 32555
rect 12894 32552 12900 32564
rect 12667 32524 12900 32552
rect 12667 32521 12679 32524
rect 12621 32515 12679 32521
rect 12894 32512 12900 32524
rect 12952 32512 12958 32564
rect 13449 32555 13507 32561
rect 13449 32521 13461 32555
rect 13495 32552 13507 32555
rect 15286 32552 15292 32564
rect 13495 32524 15292 32552
rect 13495 32521 13507 32524
rect 13449 32515 13507 32521
rect 15286 32512 15292 32524
rect 15344 32512 15350 32564
rect 19889 32555 19947 32561
rect 19889 32521 19901 32555
rect 19935 32552 19947 32555
rect 19978 32552 19984 32564
rect 19935 32524 19984 32552
rect 19935 32521 19947 32524
rect 19889 32515 19947 32521
rect 19978 32512 19984 32524
rect 20036 32512 20042 32564
rect 20714 32512 20720 32564
rect 20772 32512 20778 32564
rect 22186 32512 22192 32564
rect 22244 32512 22250 32564
rect 24854 32512 24860 32564
rect 24912 32552 24918 32564
rect 25041 32555 25099 32561
rect 25041 32552 25053 32555
rect 24912 32524 25053 32552
rect 24912 32512 24918 32524
rect 25041 32521 25053 32524
rect 25087 32521 25099 32555
rect 25041 32515 25099 32521
rect 25590 32512 25596 32564
rect 25648 32552 25654 32564
rect 26050 32552 26056 32564
rect 25648 32524 26056 32552
rect 25648 32512 25654 32524
rect 26050 32512 26056 32524
rect 26108 32552 26114 32564
rect 26513 32555 26571 32561
rect 26513 32552 26525 32555
rect 26108 32524 26525 32552
rect 26108 32512 26114 32524
rect 26513 32521 26525 32524
rect 26559 32521 26571 32555
rect 26513 32515 26571 32521
rect 27982 32512 27988 32564
rect 28040 32552 28046 32564
rect 28353 32555 28411 32561
rect 28353 32552 28365 32555
rect 28040 32524 28365 32552
rect 28040 32512 28046 32524
rect 28353 32521 28365 32524
rect 28399 32521 28411 32555
rect 28353 32515 28411 32521
rect 13814 32444 13820 32496
rect 13872 32484 13878 32496
rect 21266 32484 21272 32496
rect 13872 32456 14412 32484
rect 13872 32444 13878 32456
rect 12161 32419 12219 32425
rect 12161 32385 12173 32419
rect 12207 32416 12219 32419
rect 12802 32416 12808 32428
rect 12207 32388 12808 32416
rect 12207 32385 12219 32388
rect 12161 32379 12219 32385
rect 12802 32376 12808 32388
rect 12860 32376 12866 32428
rect 12989 32419 13047 32425
rect 12989 32385 13001 32419
rect 13035 32416 13047 32419
rect 13541 32419 13599 32425
rect 13541 32416 13553 32419
rect 13035 32388 13553 32416
rect 13035 32385 13047 32388
rect 12989 32379 13047 32385
rect 13541 32385 13553 32388
rect 13587 32385 13599 32419
rect 13541 32379 13599 32385
rect 13630 32376 13636 32428
rect 13688 32416 13694 32428
rect 13725 32419 13783 32425
rect 13725 32416 13737 32419
rect 13688 32388 13737 32416
rect 13688 32376 13694 32388
rect 13725 32385 13737 32388
rect 13771 32385 13783 32419
rect 13725 32379 13783 32385
rect 12253 32351 12311 32357
rect 12253 32317 12265 32351
rect 12299 32348 12311 32351
rect 12526 32348 12532 32360
rect 12299 32320 12532 32348
rect 12299 32317 12311 32320
rect 12253 32311 12311 32317
rect 12526 32308 12532 32320
rect 12584 32308 12590 32360
rect 13078 32308 13084 32360
rect 13136 32308 13142 32360
rect 13170 32308 13176 32360
rect 13228 32308 13234 32360
rect 13265 32351 13323 32357
rect 13265 32317 13277 32351
rect 13311 32348 13323 32351
rect 13832 32348 13860 32444
rect 13906 32376 13912 32428
rect 13964 32416 13970 32428
rect 14001 32419 14059 32425
rect 14001 32416 14013 32419
rect 13964 32388 14013 32416
rect 13964 32376 13970 32388
rect 14001 32385 14013 32388
rect 14047 32385 14059 32419
rect 14001 32379 14059 32385
rect 13311 32320 13860 32348
rect 14016 32348 14044 32379
rect 14090 32376 14096 32428
rect 14148 32376 14154 32428
rect 14182 32376 14188 32428
rect 14240 32376 14246 32428
rect 14384 32425 14412 32456
rect 20732 32456 21272 32484
rect 14369 32419 14427 32425
rect 14369 32385 14381 32419
rect 14415 32385 14427 32419
rect 14369 32379 14427 32385
rect 14645 32419 14703 32425
rect 14645 32385 14657 32419
rect 14691 32385 14703 32419
rect 14645 32379 14703 32385
rect 14660 32348 14688 32379
rect 19242 32376 19248 32428
rect 19300 32376 19306 32428
rect 20732 32425 20760 32456
rect 21266 32444 21272 32456
rect 21324 32444 21330 32496
rect 21818 32444 21824 32496
rect 21876 32484 21882 32496
rect 21876 32456 27016 32484
rect 21876 32444 21882 32456
rect 20717 32419 20775 32425
rect 20717 32385 20729 32419
rect 20763 32385 20775 32419
rect 20717 32379 20775 32385
rect 20806 32376 20812 32428
rect 20864 32376 20870 32428
rect 20990 32376 20996 32428
rect 21048 32376 21054 32428
rect 22370 32376 22376 32428
rect 22428 32376 22434 32428
rect 22462 32376 22468 32428
rect 22520 32416 22526 32428
rect 22557 32419 22615 32425
rect 22557 32416 22569 32419
rect 22520 32388 22569 32416
rect 22520 32376 22526 32388
rect 22557 32385 22569 32388
rect 22603 32385 22615 32419
rect 22557 32379 22615 32385
rect 22649 32419 22707 32425
rect 22649 32385 22661 32419
rect 22695 32416 22707 32419
rect 23290 32416 23296 32428
rect 22695 32388 23296 32416
rect 22695 32385 22707 32388
rect 22649 32379 22707 32385
rect 23290 32376 23296 32388
rect 23348 32376 23354 32428
rect 23676 32425 23704 32456
rect 23661 32419 23719 32425
rect 23661 32385 23673 32419
rect 23707 32385 23719 32419
rect 23661 32379 23719 32385
rect 23928 32419 23986 32425
rect 23928 32385 23940 32419
rect 23974 32416 23986 32419
rect 24394 32416 24400 32428
rect 23974 32388 24400 32416
rect 23974 32385 23986 32388
rect 23928 32379 23986 32385
rect 24394 32376 24400 32388
rect 24452 32376 24458 32428
rect 25148 32425 25176 32456
rect 26988 32428 27016 32456
rect 25406 32425 25412 32428
rect 25133 32419 25191 32425
rect 25133 32385 25145 32419
rect 25179 32385 25191 32419
rect 25133 32379 25191 32385
rect 25400 32379 25412 32425
rect 25406 32376 25412 32379
rect 25464 32376 25470 32428
rect 26970 32376 26976 32428
rect 27028 32376 27034 32428
rect 27062 32376 27068 32428
rect 27120 32416 27126 32428
rect 27229 32419 27287 32425
rect 27229 32416 27241 32419
rect 27120 32388 27241 32416
rect 27120 32376 27126 32388
rect 27229 32385 27241 32388
rect 27275 32385 27287 32419
rect 27229 32379 27287 32385
rect 14016 32320 14688 32348
rect 13311 32317 13323 32320
rect 13265 32311 13323 32317
rect 12986 32240 12992 32292
rect 13044 32280 13050 32292
rect 13280 32280 13308 32311
rect 14553 32283 14611 32289
rect 14553 32280 14565 32283
rect 13044 32252 13308 32280
rect 13556 32252 14565 32280
rect 13044 32240 13050 32252
rect 842 32172 848 32224
rect 900 32212 906 32224
rect 1397 32215 1455 32221
rect 1397 32212 1409 32215
rect 900 32184 1409 32212
rect 900 32172 906 32184
rect 1397 32181 1409 32184
rect 1443 32181 1455 32215
rect 1397 32175 1455 32181
rect 11974 32172 11980 32224
rect 12032 32172 12038 32224
rect 12434 32172 12440 32224
rect 12492 32212 12498 32224
rect 13556 32212 13584 32252
rect 14553 32249 14565 32252
rect 14599 32249 14611 32283
rect 14553 32243 14611 32249
rect 12492 32184 13584 32212
rect 12492 32172 12498 32184
rect 13814 32172 13820 32224
rect 13872 32212 13878 32224
rect 13909 32215 13967 32221
rect 13909 32212 13921 32215
rect 13872 32184 13921 32212
rect 13872 32172 13878 32184
rect 13909 32181 13921 32184
rect 13955 32181 13967 32215
rect 13909 32175 13967 32181
rect 13998 32172 14004 32224
rect 14056 32212 14062 32224
rect 14737 32215 14795 32221
rect 14737 32212 14749 32215
rect 14056 32184 14749 32212
rect 14056 32172 14062 32184
rect 14737 32181 14749 32184
rect 14783 32212 14795 32215
rect 17862 32212 17868 32224
rect 14783 32184 17868 32212
rect 14783 32181 14795 32184
rect 14737 32175 14795 32181
rect 17862 32172 17868 32184
rect 17920 32172 17926 32224
rect 1104 32122 28888 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 28888 32122
rect 1104 32048 28888 32070
rect 12986 31968 12992 32020
rect 13044 31968 13050 32020
rect 13078 31968 13084 32020
rect 13136 32008 13142 32020
rect 14093 32011 14151 32017
rect 14093 32008 14105 32011
rect 13136 31980 14105 32008
rect 13136 31968 13142 31980
rect 14093 31977 14105 31980
rect 14139 31977 14151 32011
rect 14093 31971 14151 31977
rect 24394 31968 24400 32020
rect 24452 31968 24458 32020
rect 24762 31968 24768 32020
rect 24820 31968 24826 32020
rect 26142 31968 26148 32020
rect 26200 32008 26206 32020
rect 26605 32011 26663 32017
rect 26605 32008 26617 32011
rect 26200 31980 26617 32008
rect 26200 31968 26206 31980
rect 26605 31977 26617 31980
rect 26651 31977 26663 32011
rect 26605 31971 26663 31977
rect 26973 32011 27031 32017
rect 26973 31977 26985 32011
rect 27019 32008 27031 32011
rect 27062 32008 27068 32020
rect 27019 31980 27068 32008
rect 27019 31977 27031 31980
rect 26973 31971 27031 31977
rect 27062 31968 27068 31980
rect 27120 31968 27126 32020
rect 11793 31943 11851 31949
rect 11793 31909 11805 31943
rect 11839 31940 11851 31943
rect 14182 31940 14188 31952
rect 11839 31912 14188 31940
rect 11839 31909 11851 31912
rect 11793 31903 11851 31909
rect 14182 31900 14188 31912
rect 14240 31940 14246 31952
rect 14240 31912 14412 31940
rect 14240 31900 14246 31912
rect 12710 31872 12716 31884
rect 11900 31844 12716 31872
rect 842 31764 848 31816
rect 900 31804 906 31816
rect 1397 31807 1455 31813
rect 1397 31804 1409 31807
rect 900 31776 1409 31804
rect 900 31764 906 31776
rect 1397 31773 1409 31776
rect 1443 31773 1455 31807
rect 1397 31767 1455 31773
rect 8846 31764 8852 31816
rect 8904 31804 8910 31816
rect 8941 31807 8999 31813
rect 8941 31804 8953 31807
rect 8904 31776 8953 31804
rect 8904 31764 8910 31776
rect 8941 31773 8953 31776
rect 8987 31773 8999 31807
rect 8941 31767 8999 31773
rect 11698 31764 11704 31816
rect 11756 31764 11762 31816
rect 11900 31813 11928 31844
rect 12710 31832 12716 31844
rect 12768 31832 12774 31884
rect 12805 31875 12863 31881
rect 12805 31841 12817 31875
rect 12851 31872 12863 31875
rect 12851 31844 13124 31872
rect 12851 31841 12863 31844
rect 12805 31835 12863 31841
rect 11885 31807 11943 31813
rect 11885 31773 11897 31807
rect 11931 31773 11943 31807
rect 11885 31767 11943 31773
rect 12529 31807 12587 31813
rect 12529 31773 12541 31807
rect 12575 31804 12587 31807
rect 12894 31804 12900 31816
rect 12575 31776 12900 31804
rect 12575 31773 12587 31776
rect 12529 31767 12587 31773
rect 12894 31764 12900 31776
rect 12952 31764 12958 31816
rect 8662 31696 8668 31748
rect 8720 31736 8726 31748
rect 9186 31739 9244 31745
rect 9186 31736 9198 31739
rect 8720 31708 9198 31736
rect 8720 31696 8726 31708
rect 9186 31705 9198 31708
rect 9232 31705 9244 31739
rect 9186 31699 9244 31705
rect 10318 31628 10324 31680
rect 10376 31628 10382 31680
rect 13096 31668 13124 31844
rect 13354 31832 13360 31884
rect 13412 31832 13418 31884
rect 13998 31872 14004 31884
rect 13832 31844 14004 31872
rect 13265 31807 13323 31813
rect 13265 31773 13277 31807
rect 13311 31804 13323 31807
rect 13832 31804 13860 31844
rect 13998 31832 14004 31844
rect 14056 31832 14062 31884
rect 14384 31813 14412 31912
rect 20898 31900 20904 31952
rect 20956 31940 20962 31952
rect 21266 31940 21272 31952
rect 20956 31912 21272 31940
rect 20956 31900 20962 31912
rect 21266 31900 21272 31912
rect 21324 31940 21330 31952
rect 24302 31940 24308 31952
rect 21324 31912 22094 31940
rect 21324 31900 21330 31912
rect 13311 31776 13860 31804
rect 13909 31807 13967 31813
rect 13311 31773 13323 31776
rect 13265 31767 13323 31773
rect 13909 31773 13921 31807
rect 13955 31804 13967 31807
rect 14277 31807 14335 31813
rect 14277 31804 14289 31807
rect 13955 31776 14289 31804
rect 13955 31773 13967 31776
rect 13909 31767 13967 31773
rect 14277 31773 14289 31776
rect 14323 31773 14335 31807
rect 14277 31767 14335 31773
rect 14369 31807 14427 31813
rect 14369 31773 14381 31807
rect 14415 31773 14427 31807
rect 14369 31767 14427 31773
rect 16298 31764 16304 31816
rect 16356 31804 16362 31816
rect 16574 31804 16580 31816
rect 16356 31776 16580 31804
rect 16356 31764 16362 31776
rect 16574 31764 16580 31776
rect 16632 31764 16638 31816
rect 22066 31804 22094 31912
rect 24044 31912 24308 31940
rect 24044 31813 24072 31912
rect 24302 31900 24308 31912
rect 24360 31940 24366 31952
rect 24360 31912 24808 31940
rect 24360 31900 24366 31912
rect 24121 31875 24179 31881
rect 24121 31841 24133 31875
rect 24167 31872 24179 31875
rect 24780 31872 24808 31912
rect 24854 31900 24860 31952
rect 24912 31940 24918 31952
rect 24912 31912 25544 31940
rect 24912 31900 24918 31912
rect 25516 31881 25544 31912
rect 28442 31900 28448 31952
rect 28500 31900 28506 31952
rect 25501 31875 25559 31881
rect 24167 31844 24624 31872
rect 24780 31844 25452 31872
rect 24167 31841 24179 31844
rect 24121 31835 24179 31841
rect 24029 31807 24087 31813
rect 24029 31804 24041 31807
rect 22066 31776 24041 31804
rect 24029 31773 24041 31776
rect 24075 31773 24087 31807
rect 24029 31767 24087 31773
rect 24210 31764 24216 31816
rect 24268 31804 24274 31816
rect 24596 31813 24624 31844
rect 24581 31807 24639 31813
rect 24268 31776 24532 31804
rect 24268 31764 24274 31776
rect 13538 31696 13544 31748
rect 13596 31696 13602 31748
rect 13725 31739 13783 31745
rect 13725 31705 13737 31739
rect 13771 31736 13783 31739
rect 13814 31736 13820 31748
rect 13771 31708 13820 31736
rect 13771 31705 13783 31708
rect 13725 31699 13783 31705
rect 13814 31696 13820 31708
rect 13872 31696 13878 31748
rect 24504 31736 24532 31776
rect 24581 31773 24593 31807
rect 24627 31773 24639 31807
rect 24581 31767 24639 31773
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 24949 31807 25007 31813
rect 24949 31804 24961 31807
rect 24903 31776 24961 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 24949 31773 24961 31776
rect 24995 31773 25007 31807
rect 25424 31804 25452 31844
rect 25501 31841 25513 31875
rect 25547 31841 25559 31875
rect 25501 31835 25559 31841
rect 26050 31832 26056 31884
rect 26108 31872 26114 31884
rect 26329 31875 26387 31881
rect 26329 31872 26341 31875
rect 26108 31844 26341 31872
rect 26108 31832 26114 31844
rect 26329 31841 26341 31844
rect 26375 31841 26387 31875
rect 26329 31835 26387 31841
rect 26510 31832 26516 31884
rect 26568 31832 26574 31884
rect 25682 31804 25688 31816
rect 25424 31776 25688 31804
rect 24949 31767 25007 31773
rect 25682 31764 25688 31776
rect 25740 31764 25746 31816
rect 26786 31764 26792 31816
rect 26844 31764 26850 31816
rect 28261 31807 28319 31813
rect 28261 31773 28273 31807
rect 28307 31804 28319 31807
rect 28350 31804 28356 31816
rect 28307 31776 28356 31804
rect 28307 31773 28319 31776
rect 28261 31767 28319 31773
rect 28350 31764 28356 31776
rect 28408 31764 28414 31816
rect 25038 31736 25044 31748
rect 24504 31708 25044 31736
rect 25038 31696 25044 31708
rect 25096 31696 25102 31748
rect 13262 31668 13268 31680
rect 13096 31640 13268 31668
rect 13262 31628 13268 31640
rect 13320 31628 13326 31680
rect 24946 31628 24952 31680
rect 25004 31668 25010 31680
rect 25777 31671 25835 31677
rect 25777 31668 25789 31671
rect 25004 31640 25789 31668
rect 25004 31628 25010 31640
rect 25777 31637 25789 31640
rect 25823 31637 25835 31671
rect 25777 31631 25835 31637
rect 1104 31578 28888 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 28888 31578
rect 1104 31504 28888 31526
rect 8662 31424 8668 31476
rect 8720 31424 8726 31476
rect 12802 31424 12808 31476
rect 12860 31464 12866 31476
rect 13541 31467 13599 31473
rect 13541 31464 13553 31467
rect 12860 31436 13553 31464
rect 12860 31424 12866 31436
rect 13541 31433 13553 31436
rect 13587 31433 13599 31467
rect 13541 31427 13599 31433
rect 25406 31424 25412 31476
rect 25464 31424 25470 31476
rect 8570 31396 8576 31408
rect 8496 31368 8576 31396
rect 5629 31331 5687 31337
rect 5629 31297 5641 31331
rect 5675 31328 5687 31331
rect 6549 31331 6607 31337
rect 6549 31328 6561 31331
rect 5675 31300 6561 31328
rect 5675 31297 5687 31300
rect 5629 31291 5687 31297
rect 6549 31297 6561 31300
rect 6595 31328 6607 31331
rect 6914 31328 6920 31340
rect 6595 31300 6920 31328
rect 6595 31297 6607 31300
rect 6549 31291 6607 31297
rect 6914 31288 6920 31300
rect 6972 31288 6978 31340
rect 8496 31337 8524 31368
rect 8570 31356 8576 31368
rect 8628 31396 8634 31408
rect 8628 31368 12204 31396
rect 8628 31356 8634 31368
rect 8481 31331 8539 31337
rect 8481 31297 8493 31331
rect 8527 31297 8539 31331
rect 8481 31291 8539 31297
rect 11698 31288 11704 31340
rect 11756 31328 11762 31340
rect 11793 31331 11851 31337
rect 11793 31328 11805 31331
rect 11756 31300 11805 31328
rect 11756 31288 11762 31300
rect 11793 31297 11805 31300
rect 11839 31297 11851 31331
rect 11793 31291 11851 31297
rect 5810 31220 5816 31272
rect 5868 31220 5874 31272
rect 6454 31220 6460 31272
rect 6512 31260 6518 31272
rect 6733 31263 6791 31269
rect 6733 31260 6745 31263
rect 6512 31232 6745 31260
rect 6512 31220 6518 31232
rect 6733 31229 6745 31232
rect 6779 31229 6791 31263
rect 6733 31223 6791 31229
rect 8297 31263 8355 31269
rect 8297 31229 8309 31263
rect 8343 31260 8355 31263
rect 8757 31263 8815 31269
rect 8757 31260 8769 31263
rect 8343 31232 8769 31260
rect 8343 31229 8355 31232
rect 8297 31223 8355 31229
rect 8757 31229 8769 31232
rect 8803 31229 8815 31263
rect 8757 31223 8815 31229
rect 9214 31220 9220 31272
rect 9272 31260 9278 31272
rect 9309 31263 9367 31269
rect 9309 31260 9321 31263
rect 9272 31232 9321 31260
rect 9272 31220 9278 31232
rect 9309 31229 9321 31232
rect 9355 31229 9367 31263
rect 11808 31260 11836 31291
rect 11882 31288 11888 31340
rect 11940 31288 11946 31340
rect 11974 31288 11980 31340
rect 12032 31288 12038 31340
rect 12176 31337 12204 31368
rect 12710 31356 12716 31408
rect 12768 31396 12774 31408
rect 13078 31396 13084 31408
rect 12768 31368 13084 31396
rect 12768 31356 12774 31368
rect 13078 31356 13084 31368
rect 13136 31396 13142 31408
rect 13357 31399 13415 31405
rect 13357 31396 13369 31399
rect 13136 31368 13369 31396
rect 13136 31356 13142 31368
rect 13357 31365 13369 31368
rect 13403 31365 13415 31399
rect 25593 31399 25651 31405
rect 25593 31396 25605 31399
rect 13357 31359 13415 31365
rect 25240 31368 25605 31396
rect 12161 31331 12219 31337
rect 12161 31297 12173 31331
rect 12207 31328 12219 31331
rect 12434 31328 12440 31340
rect 12207 31300 12440 31328
rect 12207 31297 12219 31300
rect 12161 31291 12219 31297
rect 12434 31288 12440 31300
rect 12492 31328 12498 31340
rect 12618 31328 12624 31340
rect 12492 31300 12624 31328
rect 12492 31288 12498 31300
rect 12618 31288 12624 31300
rect 12676 31328 12682 31340
rect 12805 31331 12863 31337
rect 12805 31328 12817 31331
rect 12676 31300 12817 31328
rect 12676 31288 12682 31300
rect 12805 31297 12817 31300
rect 12851 31297 12863 31331
rect 12805 31291 12863 31297
rect 12894 31288 12900 31340
rect 12952 31328 12958 31340
rect 13170 31328 13176 31340
rect 12952 31300 13176 31328
rect 12952 31288 12958 31300
rect 13170 31288 13176 31300
rect 13228 31288 13234 31340
rect 24946 31288 24952 31340
rect 25004 31288 25010 31340
rect 25038 31288 25044 31340
rect 25096 31288 25102 31340
rect 25240 31337 25268 31368
rect 25593 31365 25605 31368
rect 25639 31365 25651 31399
rect 25593 31359 25651 31365
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31297 25283 31331
rect 25225 31291 25283 31297
rect 25501 31331 25559 31337
rect 25501 31297 25513 31331
rect 25547 31297 25559 31331
rect 25501 31291 25559 31297
rect 13081 31263 13139 31269
rect 11808 31232 12434 31260
rect 9309 31223 9367 31229
rect 12406 31192 12434 31232
rect 13081 31229 13093 31263
rect 13127 31229 13139 31263
rect 25516 31260 25544 31291
rect 25682 31288 25688 31340
rect 25740 31288 25746 31340
rect 26142 31260 26148 31272
rect 25516 31232 26148 31260
rect 13081 31223 13139 31229
rect 12618 31192 12624 31204
rect 12406 31164 12624 31192
rect 12618 31152 12624 31164
rect 12676 31152 12682 31204
rect 12802 31152 12808 31204
rect 12860 31192 12866 31204
rect 13096 31192 13124 31223
rect 26142 31220 26148 31232
rect 26200 31220 26206 31272
rect 12860 31164 13124 31192
rect 12860 31152 12866 31164
rect 5442 31084 5448 31136
rect 5500 31084 5506 31136
rect 6362 31084 6368 31136
rect 6420 31084 6426 31136
rect 11514 31084 11520 31136
rect 11572 31084 11578 31136
rect 1104 31034 28888 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 28888 31034
rect 1104 30960 28888 30982
rect 6454 30880 6460 30932
rect 6512 30880 6518 30932
rect 12526 30880 12532 30932
rect 12584 30920 12590 30932
rect 12805 30923 12863 30929
rect 12805 30920 12817 30923
rect 12584 30892 12817 30920
rect 12584 30880 12590 30892
rect 12805 30889 12817 30892
rect 12851 30889 12863 30923
rect 12805 30883 12863 30889
rect 842 30744 848 30796
rect 900 30784 906 30796
rect 1397 30787 1455 30793
rect 1397 30784 1409 30787
rect 900 30756 1409 30784
rect 900 30744 906 30756
rect 1397 30753 1409 30756
rect 1443 30753 1455 30787
rect 1397 30747 1455 30753
rect 5261 30787 5319 30793
rect 5261 30753 5273 30787
rect 5307 30784 5319 30787
rect 5721 30787 5779 30793
rect 5721 30784 5733 30787
rect 5307 30756 5733 30784
rect 5307 30753 5319 30756
rect 5261 30747 5319 30753
rect 5721 30753 5733 30756
rect 5767 30753 5779 30787
rect 6914 30784 6920 30796
rect 5721 30747 5779 30753
rect 5828 30756 6920 30784
rect 2958 30676 2964 30728
rect 3016 30716 3022 30728
rect 5445 30719 5503 30725
rect 5445 30716 5457 30719
rect 3016 30688 5457 30716
rect 3016 30676 3022 30688
rect 5445 30685 5457 30688
rect 5491 30716 5503 30719
rect 5828 30716 5856 30756
rect 6914 30744 6920 30756
rect 6972 30744 6978 30796
rect 7098 30744 7104 30796
rect 7156 30784 7162 30796
rect 7193 30787 7251 30793
rect 7193 30784 7205 30787
rect 7156 30756 7205 30784
rect 7156 30744 7162 30756
rect 7193 30753 7205 30756
rect 7239 30753 7251 30787
rect 7193 30747 7251 30753
rect 15654 30744 15660 30796
rect 15712 30744 15718 30796
rect 5491 30688 5856 30716
rect 6365 30719 6423 30725
rect 5491 30685 5503 30688
rect 5445 30679 5503 30685
rect 6365 30685 6377 30719
rect 6411 30716 6423 30719
rect 6730 30716 6736 30728
rect 6411 30688 6736 30716
rect 6411 30685 6423 30688
rect 6365 30679 6423 30685
rect 6730 30676 6736 30688
rect 6788 30716 6794 30728
rect 7469 30719 7527 30725
rect 7469 30716 7481 30719
rect 6788 30688 6914 30716
rect 6788 30676 6794 30688
rect 6886 30648 6914 30688
rect 7116 30688 7481 30716
rect 7116 30648 7144 30688
rect 7469 30685 7481 30688
rect 7515 30685 7527 30719
rect 7469 30679 7527 30685
rect 9582 30676 9588 30728
rect 9640 30716 9646 30728
rect 11514 30725 11520 30728
rect 11241 30719 11299 30725
rect 11241 30716 11253 30719
rect 9640 30688 11253 30716
rect 9640 30676 9646 30688
rect 11241 30685 11253 30688
rect 11287 30685 11299 30719
rect 11508 30716 11520 30725
rect 11475 30688 11520 30716
rect 11241 30679 11299 30685
rect 11508 30679 11520 30688
rect 11514 30676 11520 30679
rect 11572 30676 11578 30728
rect 12710 30676 12716 30728
rect 12768 30676 12774 30728
rect 12894 30676 12900 30728
rect 12952 30676 12958 30728
rect 15562 30676 15568 30728
rect 15620 30676 15626 30728
rect 6886 30620 7144 30648
rect 7561 30651 7619 30657
rect 7561 30617 7573 30651
rect 7607 30648 7619 30651
rect 9214 30648 9220 30660
rect 7607 30620 9220 30648
rect 7607 30617 7619 30620
rect 7561 30611 7619 30617
rect 9214 30608 9220 30620
rect 9272 30608 9278 30660
rect 5629 30583 5687 30589
rect 5629 30549 5641 30583
rect 5675 30580 5687 30583
rect 6638 30580 6644 30592
rect 5675 30552 6644 30580
rect 5675 30549 5687 30552
rect 5629 30543 5687 30549
rect 6638 30540 6644 30552
rect 6696 30540 6702 30592
rect 6914 30540 6920 30592
rect 6972 30580 6978 30592
rect 7377 30583 7435 30589
rect 7377 30580 7389 30583
rect 6972 30552 7389 30580
rect 6972 30540 6978 30552
rect 7377 30549 7389 30552
rect 7423 30549 7435 30583
rect 7377 30543 7435 30549
rect 7745 30583 7803 30589
rect 7745 30549 7757 30583
rect 7791 30580 7803 30583
rect 8938 30580 8944 30592
rect 7791 30552 8944 30580
rect 7791 30549 7803 30552
rect 7745 30543 7803 30549
rect 8938 30540 8944 30552
rect 8996 30540 9002 30592
rect 12618 30540 12624 30592
rect 12676 30580 12682 30592
rect 13814 30580 13820 30592
rect 12676 30552 13820 30580
rect 12676 30540 12682 30552
rect 13814 30540 13820 30552
rect 13872 30580 13878 30592
rect 15102 30580 15108 30592
rect 13872 30552 15108 30580
rect 13872 30540 13878 30552
rect 15102 30540 15108 30552
rect 15160 30540 15166 30592
rect 15930 30540 15936 30592
rect 15988 30540 15994 30592
rect 1104 30490 28888 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 28888 30490
rect 1104 30416 28888 30438
rect 11882 30336 11888 30388
rect 11940 30376 11946 30388
rect 13630 30376 13636 30388
rect 11940 30348 13636 30376
rect 11940 30336 11946 30348
rect 13630 30336 13636 30348
rect 13688 30336 13694 30388
rect 6638 30317 6644 30320
rect 6632 30308 6644 30317
rect 4816 30280 6408 30308
rect 6599 30280 6644 30308
rect 4706 30132 4712 30184
rect 4764 30172 4770 30184
rect 4816 30181 4844 30280
rect 5068 30243 5126 30249
rect 5068 30209 5080 30243
rect 5114 30240 5126 30243
rect 5442 30240 5448 30252
rect 5114 30212 5448 30240
rect 5114 30209 5126 30212
rect 5068 30203 5126 30209
rect 5442 30200 5448 30212
rect 5500 30200 5506 30252
rect 6380 30249 6408 30280
rect 6632 30271 6644 30280
rect 6638 30268 6644 30271
rect 6696 30268 6702 30320
rect 8846 30268 8852 30320
rect 8904 30308 8910 30320
rect 9582 30308 9588 30320
rect 8904 30280 9588 30308
rect 8904 30268 8910 30280
rect 9582 30268 9588 30280
rect 9640 30308 9646 30320
rect 15749 30311 15807 30317
rect 9640 30280 10272 30308
rect 9640 30268 9646 30280
rect 6365 30243 6423 30249
rect 6365 30209 6377 30243
rect 6411 30209 6423 30243
rect 6365 30203 6423 30209
rect 7006 30200 7012 30252
rect 7064 30240 7070 30252
rect 7374 30240 7380 30252
rect 7064 30212 7380 30240
rect 7064 30200 7070 30212
rect 7374 30200 7380 30212
rect 7432 30240 7438 30252
rect 10244 30249 10272 30280
rect 15749 30277 15761 30311
rect 15795 30308 15807 30311
rect 15930 30308 15936 30320
rect 15795 30280 15936 30308
rect 15795 30277 15807 30280
rect 15749 30271 15807 30277
rect 15930 30268 15936 30280
rect 15988 30268 15994 30320
rect 9973 30243 10031 30249
rect 7432 30212 9260 30240
rect 7432 30200 7438 30212
rect 4801 30175 4859 30181
rect 4801 30172 4813 30175
rect 4764 30144 4813 30172
rect 4764 30132 4770 30144
rect 4801 30141 4813 30144
rect 4847 30141 4859 30175
rect 8389 30175 8447 30181
rect 8389 30172 8401 30175
rect 4801 30135 4859 30141
rect 7760 30144 8401 30172
rect 7760 30116 7788 30144
rect 8389 30141 8401 30144
rect 8435 30141 8447 30175
rect 8389 30135 8447 30141
rect 7742 30064 7748 30116
rect 7800 30064 7806 30116
rect 9232 30104 9260 30212
rect 9973 30209 9985 30243
rect 10019 30240 10031 30243
rect 10229 30243 10287 30249
rect 10019 30212 10180 30240
rect 10019 30209 10031 30212
rect 9973 30203 10031 30209
rect 10152 30172 10180 30212
rect 10229 30209 10241 30243
rect 10275 30209 10287 30243
rect 10229 30203 10287 30209
rect 10505 30243 10563 30249
rect 10505 30209 10517 30243
rect 10551 30209 10563 30243
rect 10505 30203 10563 30209
rect 10321 30175 10379 30181
rect 10321 30172 10333 30175
rect 10152 30144 10333 30172
rect 10321 30141 10333 30144
rect 10367 30141 10379 30175
rect 10321 30135 10379 30141
rect 9232 30076 9352 30104
rect 6181 30039 6239 30045
rect 6181 30005 6193 30039
rect 6227 30036 6239 30039
rect 7098 30036 7104 30048
rect 6227 30008 7104 30036
rect 6227 30005 6239 30008
rect 6181 29999 6239 30005
rect 7098 29996 7104 30008
rect 7156 29996 7162 30048
rect 7282 29996 7288 30048
rect 7340 30036 7346 30048
rect 7837 30039 7895 30045
rect 7837 30036 7849 30039
rect 7340 30008 7849 30036
rect 7340 29996 7346 30008
rect 7837 30005 7849 30008
rect 7883 30005 7895 30039
rect 7837 29999 7895 30005
rect 8849 30039 8907 30045
rect 8849 30005 8861 30039
rect 8895 30036 8907 30039
rect 9214 30036 9220 30048
rect 8895 30008 9220 30036
rect 8895 30005 8907 30008
rect 8849 29999 8907 30005
rect 9214 29996 9220 30008
rect 9272 29996 9278 30048
rect 9324 30036 9352 30076
rect 10520 30036 10548 30203
rect 15286 30200 15292 30252
rect 15344 30200 15350 30252
rect 15841 30243 15899 30249
rect 15841 30209 15853 30243
rect 15887 30240 15899 30243
rect 16298 30240 16304 30252
rect 15887 30212 16304 30240
rect 15887 30209 15899 30212
rect 15841 30203 15899 30209
rect 16298 30200 16304 30212
rect 16356 30200 16362 30252
rect 16390 30200 16396 30252
rect 16448 30240 16454 30252
rect 16485 30243 16543 30249
rect 16485 30240 16497 30243
rect 16448 30212 16497 30240
rect 16448 30200 16454 30212
rect 16485 30209 16497 30212
rect 16531 30209 16543 30243
rect 16485 30203 16543 30209
rect 26970 30200 26976 30252
rect 27028 30200 27034 30252
rect 27062 30200 27068 30252
rect 27120 30240 27126 30252
rect 27229 30243 27287 30249
rect 27229 30240 27241 30243
rect 27120 30212 27241 30240
rect 27120 30200 27126 30212
rect 27229 30209 27241 30212
rect 27275 30209 27287 30243
rect 27229 30203 27287 30209
rect 10686 30132 10692 30184
rect 10744 30132 10750 30184
rect 12618 30132 12624 30184
rect 12676 30172 12682 30184
rect 13538 30172 13544 30184
rect 12676 30144 13544 30172
rect 12676 30132 12682 30144
rect 13538 30132 13544 30144
rect 13596 30172 13602 30184
rect 15197 30175 15255 30181
rect 15197 30172 15209 30175
rect 13596 30144 15209 30172
rect 13596 30132 13602 30144
rect 15197 30141 15209 30144
rect 15243 30141 15255 30175
rect 15197 30135 15255 30141
rect 15654 30132 15660 30184
rect 15712 30132 15718 30184
rect 16117 30175 16175 30181
rect 16117 30141 16129 30175
rect 16163 30172 16175 30175
rect 19334 30172 19340 30184
rect 16163 30144 19340 30172
rect 16163 30141 16175 30144
rect 16117 30135 16175 30141
rect 19334 30132 19340 30144
rect 19392 30132 19398 30184
rect 16025 30107 16083 30113
rect 16025 30073 16037 30107
rect 16071 30104 16083 30107
rect 16301 30107 16359 30113
rect 16301 30104 16313 30107
rect 16071 30076 16313 30104
rect 16071 30073 16083 30076
rect 16025 30067 16083 30073
rect 16301 30073 16313 30076
rect 16347 30073 16359 30107
rect 16301 30067 16359 30073
rect 28350 30064 28356 30116
rect 28408 30064 28414 30116
rect 11330 30036 11336 30048
rect 9324 30008 11336 30036
rect 11330 29996 11336 30008
rect 11388 29996 11394 30048
rect 16206 29996 16212 30048
rect 16264 29996 16270 30048
rect 1104 29946 28888 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 28888 29946
rect 1104 29872 28888 29894
rect 5261 29835 5319 29841
rect 5261 29801 5273 29835
rect 5307 29832 5319 29835
rect 6822 29832 6828 29844
rect 5307 29804 6828 29832
rect 5307 29801 5319 29804
rect 5261 29795 5319 29801
rect 6822 29792 6828 29804
rect 6880 29792 6886 29844
rect 7742 29832 7748 29844
rect 6932 29804 7748 29832
rect 1581 29767 1639 29773
rect 1581 29733 1593 29767
rect 1627 29733 1639 29767
rect 1581 29727 1639 29733
rect 1596 29696 1624 29727
rect 6730 29724 6736 29776
rect 6788 29724 6794 29776
rect 6932 29705 6960 29804
rect 7742 29792 7748 29804
rect 7800 29792 7806 29844
rect 11330 29792 11336 29844
rect 11388 29792 11394 29844
rect 8757 29767 8815 29773
rect 8757 29733 8769 29767
rect 8803 29764 8815 29767
rect 8803 29736 9352 29764
rect 8803 29733 8815 29736
rect 8757 29727 8815 29733
rect 6917 29699 6975 29705
rect 1596 29668 3096 29696
rect 842 29588 848 29640
rect 900 29628 906 29640
rect 1397 29631 1455 29637
rect 1397 29628 1409 29631
rect 900 29600 1409 29628
rect 900 29588 906 29600
rect 1397 29597 1409 29600
rect 1443 29597 1455 29631
rect 1397 29591 1455 29597
rect 2958 29588 2964 29640
rect 3016 29588 3022 29640
rect 3068 29637 3096 29668
rect 6917 29665 6929 29699
rect 6963 29665 6975 29699
rect 7377 29699 7435 29705
rect 7377 29696 7389 29699
rect 6917 29659 6975 29665
rect 7024 29668 7389 29696
rect 3053 29631 3111 29637
rect 3053 29597 3065 29631
rect 3099 29597 3111 29631
rect 3053 29591 3111 29597
rect 3881 29631 3939 29637
rect 3881 29597 3893 29631
rect 3927 29628 3939 29631
rect 4706 29628 4712 29640
rect 3927 29600 4712 29628
rect 3927 29597 3939 29600
rect 3881 29591 3939 29597
rect 4706 29588 4712 29600
rect 4764 29628 4770 29640
rect 5353 29631 5411 29637
rect 5353 29628 5365 29631
rect 4764 29600 5365 29628
rect 4764 29588 4770 29600
rect 5353 29597 5365 29600
rect 5399 29628 5411 29631
rect 7024 29628 7052 29668
rect 7377 29665 7389 29668
rect 7423 29665 7435 29699
rect 7377 29659 7435 29665
rect 5399 29600 7052 29628
rect 5399 29597 5411 29600
rect 5353 29591 5411 29597
rect 7098 29588 7104 29640
rect 7156 29588 7162 29640
rect 7392 29628 7420 29659
rect 8938 29656 8944 29708
rect 8996 29656 9002 29708
rect 9324 29705 9352 29736
rect 9309 29699 9367 29705
rect 9309 29665 9321 29699
rect 9355 29696 9367 29699
rect 10229 29699 10287 29705
rect 10229 29696 10241 29699
rect 9355 29668 10241 29696
rect 9355 29665 9367 29668
rect 9309 29659 9367 29665
rect 10229 29665 10241 29668
rect 10275 29696 10287 29699
rect 10594 29696 10600 29708
rect 10275 29668 10600 29696
rect 10275 29665 10287 29668
rect 10229 29659 10287 29665
rect 10594 29656 10600 29668
rect 10652 29656 10658 29708
rect 17037 29699 17095 29705
rect 17037 29665 17049 29699
rect 17083 29696 17095 29699
rect 17770 29696 17776 29708
rect 17083 29668 17776 29696
rect 17083 29665 17095 29668
rect 17037 29659 17095 29665
rect 17770 29656 17776 29668
rect 17828 29656 17834 29708
rect 8846 29628 8852 29640
rect 7392 29600 8852 29628
rect 8846 29588 8852 29600
rect 8904 29588 8910 29640
rect 9401 29631 9459 29637
rect 9401 29597 9413 29631
rect 9447 29628 9459 29631
rect 9490 29628 9496 29640
rect 9447 29600 9496 29628
rect 9447 29597 9459 29600
rect 9401 29591 9459 29597
rect 9490 29588 9496 29600
rect 9548 29588 9554 29640
rect 10410 29588 10416 29640
rect 10468 29588 10474 29640
rect 11241 29631 11299 29637
rect 11241 29597 11253 29631
rect 11287 29628 11299 29631
rect 12342 29628 12348 29640
rect 11287 29600 12348 29628
rect 11287 29597 11299 29600
rect 11241 29591 11299 29597
rect 12342 29588 12348 29600
rect 12400 29588 12406 29640
rect 16206 29588 16212 29640
rect 16264 29628 16270 29640
rect 16770 29631 16828 29637
rect 16770 29628 16782 29631
rect 16264 29600 16782 29628
rect 16264 29588 16270 29600
rect 16770 29597 16782 29600
rect 16816 29597 16828 29631
rect 16770 29591 16828 29597
rect 3237 29563 3295 29569
rect 3237 29529 3249 29563
rect 3283 29560 3295 29563
rect 4126 29563 4184 29569
rect 4126 29560 4138 29563
rect 3283 29532 4138 29560
rect 3283 29529 3295 29532
rect 3237 29523 3295 29529
rect 4126 29529 4138 29532
rect 4172 29529 4184 29563
rect 4126 29523 4184 29529
rect 5620 29563 5678 29569
rect 5620 29529 5632 29563
rect 5666 29560 5678 29563
rect 6362 29560 6368 29572
rect 5666 29532 6368 29560
rect 5666 29529 5678 29532
rect 5620 29523 5678 29529
rect 6362 29520 6368 29532
rect 6420 29520 6426 29572
rect 6730 29520 6736 29572
rect 6788 29560 6794 29572
rect 7650 29569 7656 29572
rect 6825 29563 6883 29569
rect 6825 29560 6837 29563
rect 6788 29532 6837 29560
rect 6788 29520 6794 29532
rect 6825 29529 6837 29532
rect 6871 29529 6883 29563
rect 6825 29523 6883 29529
rect 7633 29563 7656 29569
rect 7633 29529 7645 29563
rect 7708 29560 7714 29572
rect 9033 29563 9091 29569
rect 9033 29560 9045 29563
rect 7708 29532 9045 29560
rect 7633 29523 7656 29529
rect 7650 29520 7656 29523
rect 7708 29520 7714 29532
rect 9033 29529 9045 29532
rect 9079 29529 9091 29563
rect 10318 29560 10324 29572
rect 9033 29523 9091 29529
rect 9232 29532 10324 29560
rect 7285 29495 7343 29501
rect 7285 29461 7297 29495
rect 7331 29492 7343 29495
rect 8662 29492 8668 29504
rect 7331 29464 8668 29492
rect 7331 29461 7343 29464
rect 7285 29455 7343 29461
rect 8662 29452 8668 29464
rect 8720 29452 8726 29504
rect 9232 29501 9260 29532
rect 10318 29520 10324 29532
rect 10376 29520 10382 29572
rect 9217 29495 9275 29501
rect 9217 29461 9229 29495
rect 9263 29461 9275 29495
rect 9217 29455 9275 29461
rect 9398 29452 9404 29504
rect 9456 29492 9462 29504
rect 9585 29495 9643 29501
rect 9585 29492 9597 29495
rect 9456 29464 9597 29492
rect 9456 29452 9462 29464
rect 9585 29461 9597 29464
rect 9631 29461 9643 29495
rect 9585 29455 9643 29461
rect 9674 29452 9680 29504
rect 9732 29452 9738 29504
rect 10686 29452 10692 29504
rect 10744 29492 10750 29504
rect 11057 29495 11115 29501
rect 11057 29492 11069 29495
rect 10744 29464 11069 29492
rect 10744 29452 10750 29464
rect 11057 29461 11069 29464
rect 11103 29461 11115 29495
rect 11057 29455 11115 29461
rect 15286 29452 15292 29504
rect 15344 29492 15350 29504
rect 15657 29495 15715 29501
rect 15657 29492 15669 29495
rect 15344 29464 15669 29492
rect 15344 29452 15350 29464
rect 15657 29461 15669 29464
rect 15703 29492 15715 29495
rect 16298 29492 16304 29504
rect 15703 29464 16304 29492
rect 15703 29461 15715 29464
rect 15657 29455 15715 29461
rect 16298 29452 16304 29464
rect 16356 29452 16362 29504
rect 1104 29402 28888 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 28888 29402
rect 1104 29328 28888 29350
rect 5537 29291 5595 29297
rect 5537 29257 5549 29291
rect 5583 29288 5595 29291
rect 5810 29288 5816 29300
rect 5583 29260 5816 29288
rect 5583 29257 5595 29260
rect 5537 29251 5595 29257
rect 5810 29248 5816 29260
rect 5868 29248 5874 29300
rect 7561 29291 7619 29297
rect 7561 29257 7573 29291
rect 7607 29288 7619 29291
rect 7650 29288 7656 29300
rect 7607 29260 7656 29288
rect 7607 29257 7619 29260
rect 7561 29251 7619 29257
rect 7650 29248 7656 29260
rect 7708 29248 7714 29300
rect 9674 29288 9680 29300
rect 8588 29260 9680 29288
rect 8588 29220 8616 29260
rect 9674 29248 9680 29260
rect 9732 29248 9738 29300
rect 10229 29291 10287 29297
rect 10229 29257 10241 29291
rect 10275 29288 10287 29291
rect 10410 29288 10416 29300
rect 10275 29260 10416 29288
rect 10275 29257 10287 29260
rect 10229 29251 10287 29257
rect 10410 29248 10416 29260
rect 10468 29248 10474 29300
rect 8496 29192 8616 29220
rect 8757 29223 8815 29229
rect 6181 29155 6239 29161
rect 6181 29121 6193 29155
rect 6227 29152 6239 29155
rect 6914 29152 6920 29164
rect 6227 29124 6920 29152
rect 6227 29121 6239 29124
rect 6181 29115 6239 29121
rect 6914 29112 6920 29124
rect 6972 29112 6978 29164
rect 7282 29112 7288 29164
rect 7340 29112 7346 29164
rect 7374 29112 7380 29164
rect 7432 29112 7438 29164
rect 8496 29161 8524 29192
rect 8757 29189 8769 29223
rect 8803 29220 8815 29223
rect 9094 29223 9152 29229
rect 9094 29220 9106 29223
rect 8803 29192 9106 29220
rect 8803 29189 8815 29192
rect 8757 29183 8815 29189
rect 9094 29189 9106 29192
rect 9140 29189 9152 29223
rect 9094 29183 9152 29189
rect 9214 29180 9220 29232
rect 9272 29220 9278 29232
rect 9272 29192 10548 29220
rect 9272 29180 9278 29192
rect 8481 29155 8539 29161
rect 8481 29121 8493 29155
rect 8527 29121 8539 29155
rect 8481 29115 8539 29121
rect 8570 29112 8576 29164
rect 8628 29112 8634 29164
rect 8846 29112 8852 29164
rect 8904 29112 8910 29164
rect 10520 29161 10548 29192
rect 10321 29155 10379 29161
rect 10321 29152 10333 29155
rect 8956 29124 10333 29152
rect 8662 29044 8668 29096
rect 8720 29084 8726 29096
rect 8956 29084 8984 29124
rect 10321 29121 10333 29124
rect 10367 29121 10379 29155
rect 10321 29115 10379 29121
rect 10505 29155 10563 29161
rect 10505 29121 10517 29155
rect 10551 29121 10563 29155
rect 10505 29115 10563 29121
rect 10594 29112 10600 29164
rect 10652 29112 10658 29164
rect 15102 29112 15108 29164
rect 15160 29112 15166 29164
rect 18322 29112 18328 29164
rect 18380 29112 18386 29164
rect 18414 29112 18420 29164
rect 18472 29112 18478 29164
rect 18601 29155 18659 29161
rect 18601 29121 18613 29155
rect 18647 29152 18659 29155
rect 19334 29152 19340 29164
rect 18647 29124 19340 29152
rect 18647 29121 18659 29124
rect 18601 29115 18659 29121
rect 19334 29112 19340 29124
rect 19392 29152 19398 29164
rect 19978 29152 19984 29164
rect 19392 29124 19984 29152
rect 19392 29112 19398 29124
rect 19978 29112 19984 29124
rect 20036 29112 20042 29164
rect 8720 29056 8984 29084
rect 8720 29044 8726 29056
rect 842 28976 848 29028
rect 900 29016 906 29028
rect 1397 29019 1455 29025
rect 1397 29016 1409 29019
rect 900 28988 1409 29016
rect 900 28976 906 28988
rect 1397 28985 1409 28988
rect 1443 28985 1455 29019
rect 1397 28979 1455 28985
rect 15197 29019 15255 29025
rect 15197 28985 15209 29019
rect 15243 29016 15255 29019
rect 17494 29016 17500 29028
rect 15243 28988 17500 29016
rect 15243 28985 15255 28988
rect 15197 28979 15255 28985
rect 17494 28976 17500 28988
rect 17552 28976 17558 29028
rect 18601 29019 18659 29025
rect 18601 28985 18613 29019
rect 18647 29016 18659 29019
rect 27062 29016 27068 29028
rect 18647 28988 27068 29016
rect 18647 28985 18659 28988
rect 18601 28979 18659 28985
rect 27062 28976 27068 28988
rect 27120 28976 27126 29028
rect 10318 28908 10324 28960
rect 10376 28908 10382 28960
rect 10778 28908 10784 28960
rect 10836 28908 10842 28960
rect 1104 28858 28888 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 28888 28858
rect 1104 28784 28888 28806
rect 18414 28704 18420 28756
rect 18472 28704 18478 28756
rect 21177 28679 21235 28685
rect 21177 28645 21189 28679
rect 21223 28676 21235 28679
rect 22370 28676 22376 28688
rect 21223 28648 22376 28676
rect 21223 28645 21235 28648
rect 21177 28639 21235 28645
rect 22370 28636 22376 28648
rect 22428 28636 22434 28688
rect 17586 28568 17592 28620
rect 17644 28608 17650 28620
rect 18049 28611 18107 28617
rect 17644 28580 18000 28608
rect 17644 28568 17650 28580
rect 9125 28543 9183 28549
rect 9125 28509 9137 28543
rect 9171 28540 9183 28543
rect 9398 28540 9404 28552
rect 9171 28512 9404 28540
rect 9171 28509 9183 28512
rect 9125 28503 9183 28509
rect 9398 28500 9404 28512
rect 9456 28500 9462 28552
rect 9490 28500 9496 28552
rect 9548 28500 9554 28552
rect 17773 28543 17831 28549
rect 17773 28509 17785 28543
rect 17819 28509 17831 28543
rect 17773 28503 17831 28509
rect 9217 28475 9275 28481
rect 9217 28441 9229 28475
rect 9263 28441 9275 28475
rect 9217 28435 9275 28441
rect 9309 28475 9367 28481
rect 9309 28441 9321 28475
rect 9355 28472 9367 28475
rect 10778 28472 10784 28484
rect 9355 28444 10784 28472
rect 9355 28441 9367 28444
rect 9309 28435 9367 28441
rect 8938 28364 8944 28416
rect 8996 28364 9002 28416
rect 9232 28404 9260 28435
rect 10778 28432 10784 28444
rect 10836 28432 10842 28484
rect 16298 28432 16304 28484
rect 16356 28472 16362 28484
rect 17788 28472 17816 28503
rect 17862 28500 17868 28552
rect 17920 28500 17926 28552
rect 17972 28540 18000 28580
rect 18049 28577 18061 28611
rect 18095 28608 18107 28611
rect 19426 28608 19432 28620
rect 18095 28580 19432 28608
rect 18095 28577 18107 28580
rect 18049 28571 18107 28577
rect 19426 28568 19432 28580
rect 19484 28568 19490 28620
rect 18141 28543 18199 28549
rect 18141 28540 18153 28543
rect 17972 28512 18153 28540
rect 18141 28509 18153 28512
rect 18187 28509 18199 28543
rect 18141 28503 18199 28509
rect 18230 28500 18236 28552
rect 18288 28500 18294 28552
rect 18326 28543 18384 28549
rect 18326 28509 18338 28543
rect 18372 28509 18384 28543
rect 18326 28503 18384 28509
rect 17954 28472 17960 28484
rect 16356 28444 17724 28472
rect 17788 28444 17960 28472
rect 16356 28432 16362 28444
rect 10686 28404 10692 28416
rect 9232 28376 10692 28404
rect 10686 28364 10692 28376
rect 10744 28364 10750 28416
rect 17586 28364 17592 28416
rect 17644 28364 17650 28416
rect 17696 28404 17724 28444
rect 17954 28432 17960 28444
rect 18012 28432 18018 28484
rect 18340 28404 18368 28503
rect 19794 28500 19800 28552
rect 19852 28500 19858 28552
rect 19978 28500 19984 28552
rect 20036 28500 20042 28552
rect 20898 28500 20904 28552
rect 20956 28500 20962 28552
rect 21177 28543 21235 28549
rect 21177 28509 21189 28543
rect 21223 28540 21235 28543
rect 21266 28540 21272 28552
rect 21223 28512 21272 28540
rect 21223 28509 21235 28512
rect 21177 28503 21235 28509
rect 19996 28472 20024 28500
rect 20254 28472 20260 28484
rect 19996 28444 20260 28472
rect 20254 28432 20260 28444
rect 20312 28472 20318 28484
rect 21192 28472 21220 28503
rect 21266 28500 21272 28512
rect 21324 28500 21330 28552
rect 20312 28444 21220 28472
rect 20312 28432 20318 28444
rect 17696 28376 18368 28404
rect 19334 28364 19340 28416
rect 19392 28404 19398 28416
rect 19889 28407 19947 28413
rect 19889 28404 19901 28407
rect 19392 28376 19901 28404
rect 19392 28364 19398 28376
rect 19889 28373 19901 28376
rect 19935 28373 19947 28407
rect 19889 28367 19947 28373
rect 20806 28364 20812 28416
rect 20864 28404 20870 28416
rect 20993 28407 21051 28413
rect 20993 28404 21005 28407
rect 20864 28376 21005 28404
rect 20864 28364 20870 28376
rect 20993 28373 21005 28376
rect 21039 28373 21051 28407
rect 20993 28367 21051 28373
rect 1104 28314 28888 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 28888 28314
rect 1104 28240 28888 28262
rect 18141 28203 18199 28209
rect 18141 28169 18153 28203
rect 18187 28200 18199 28203
rect 18322 28200 18328 28212
rect 18187 28172 18328 28200
rect 18187 28169 18199 28172
rect 18141 28163 18199 28169
rect 18322 28160 18328 28172
rect 18380 28160 18386 28212
rect 19426 28160 19432 28212
rect 19484 28160 19490 28212
rect 17678 28092 17684 28144
rect 17736 28132 17742 28144
rect 17865 28135 17923 28141
rect 17865 28132 17877 28135
rect 17736 28104 17877 28132
rect 17736 28092 17742 28104
rect 17865 28101 17877 28104
rect 17911 28101 17923 28135
rect 17865 28095 17923 28101
rect 17126 28024 17132 28076
rect 17184 28064 17190 28076
rect 17497 28067 17555 28073
rect 17497 28064 17509 28067
rect 17184 28036 17509 28064
rect 17184 28024 17190 28036
rect 17497 28033 17509 28036
rect 17543 28033 17555 28067
rect 17497 28027 17555 28033
rect 17586 28024 17592 28076
rect 17644 28064 17650 28076
rect 17773 28067 17831 28073
rect 17644 28036 17689 28064
rect 17644 28024 17650 28036
rect 17773 28033 17785 28067
rect 17819 28033 17831 28067
rect 17773 28027 17831 28033
rect 18003 28067 18061 28073
rect 18003 28033 18015 28067
rect 18049 28064 18061 28067
rect 19444 28064 19472 28160
rect 20564 28135 20622 28141
rect 20564 28101 20576 28135
rect 20610 28132 20622 28135
rect 22002 28132 22008 28144
rect 20610 28104 22008 28132
rect 20610 28101 20622 28104
rect 20564 28095 20622 28101
rect 22002 28092 22008 28104
rect 22060 28092 22066 28144
rect 19610 28064 19616 28076
rect 18049 28036 19616 28064
rect 18049 28033 18061 28036
rect 18003 28027 18061 28033
rect 17788 27996 17816 28027
rect 19610 28024 19616 28036
rect 19668 28064 19674 28076
rect 20809 28067 20867 28073
rect 19668 28036 20760 28064
rect 19668 28024 19674 28036
rect 18138 27996 18144 28008
rect 17788 27968 18144 27996
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 20732 27996 20760 28036
rect 20809 28033 20821 28067
rect 20855 28064 20867 28067
rect 21174 28064 21180 28076
rect 20855 28036 21180 28064
rect 20855 28033 20867 28036
rect 20809 28027 20867 28033
rect 21174 28024 21180 28036
rect 21232 28024 21238 28076
rect 20901 27999 20959 28005
rect 20901 27996 20913 27999
rect 20732 27968 20913 27996
rect 20901 27965 20913 27968
rect 20947 27965 20959 27999
rect 20901 27959 20959 27965
rect 28534 27888 28540 27940
rect 28592 27888 28598 27940
rect 21542 27820 21548 27872
rect 21600 27820 21606 27872
rect 1104 27770 28888 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 28888 27770
rect 1104 27696 28888 27718
rect 18230 27656 18236 27668
rect 18064 27628 18236 27656
rect 16758 27548 16764 27600
rect 16816 27588 16822 27600
rect 16945 27591 17003 27597
rect 16945 27588 16957 27591
rect 16816 27560 16957 27588
rect 16816 27548 16822 27560
rect 16945 27557 16957 27560
rect 16991 27588 17003 27591
rect 18064 27588 18092 27628
rect 18230 27616 18236 27628
rect 18288 27616 18294 27668
rect 19702 27616 19708 27668
rect 19760 27656 19766 27668
rect 19760 27628 20392 27656
rect 19760 27616 19766 27628
rect 16991 27560 18092 27588
rect 16991 27557 17003 27560
rect 16945 27551 17003 27557
rect 18138 27548 18144 27600
rect 18196 27548 18202 27600
rect 19334 27548 19340 27600
rect 19392 27548 19398 27600
rect 19352 27520 19380 27548
rect 18800 27492 19380 27520
rect 20364 27520 20392 27628
rect 20898 27616 20904 27668
rect 20956 27656 20962 27668
rect 20956 27628 22232 27656
rect 20956 27616 20962 27628
rect 22204 27597 22232 27628
rect 21453 27591 21511 27597
rect 21453 27557 21465 27591
rect 21499 27588 21511 27591
rect 22189 27591 22247 27597
rect 21499 27560 22140 27588
rect 21499 27557 21511 27560
rect 21453 27551 21511 27557
rect 20364 27492 20944 27520
rect 13446 27412 13452 27464
rect 13504 27412 13510 27464
rect 13630 27412 13636 27464
rect 13688 27412 13694 27464
rect 17586 27412 17592 27464
rect 17644 27412 17650 27464
rect 17862 27412 17868 27464
rect 17920 27412 17926 27464
rect 17954 27412 17960 27464
rect 18012 27412 18018 27464
rect 18800 27461 18828 27492
rect 18785 27455 18843 27461
rect 18785 27421 18797 27455
rect 18831 27421 18843 27455
rect 18785 27415 18843 27421
rect 18966 27412 18972 27464
rect 19024 27412 19030 27464
rect 19058 27412 19064 27464
rect 19116 27412 19122 27464
rect 19337 27455 19395 27461
rect 19337 27421 19349 27455
rect 19383 27452 19395 27455
rect 19383 27424 20668 27452
rect 19383 27421 19395 27424
rect 19337 27415 19395 27421
rect 16298 27344 16304 27396
rect 16356 27384 16362 27396
rect 16669 27387 16727 27393
rect 16669 27384 16681 27387
rect 16356 27356 16681 27384
rect 16356 27344 16362 27356
rect 16669 27353 16681 27356
rect 16715 27353 16727 27387
rect 16669 27347 16727 27353
rect 17678 27344 17684 27396
rect 17736 27384 17742 27396
rect 17773 27387 17831 27393
rect 17773 27384 17785 27387
rect 17736 27356 17785 27384
rect 17736 27344 17742 27356
rect 17773 27353 17785 27356
rect 17819 27353 17831 27387
rect 17773 27347 17831 27353
rect 18601 27387 18659 27393
rect 18601 27353 18613 27387
rect 18647 27384 18659 27387
rect 19582 27387 19640 27393
rect 19582 27384 19594 27387
rect 18647 27356 19594 27384
rect 18647 27353 18659 27356
rect 18601 27347 18659 27353
rect 19582 27353 19594 27356
rect 19628 27353 19640 27387
rect 20640 27384 20668 27424
rect 20806 27412 20812 27464
rect 20864 27412 20870 27464
rect 20916 27452 20944 27492
rect 21542 27480 21548 27532
rect 21600 27480 21606 27532
rect 22002 27480 22008 27532
rect 22060 27480 22066 27532
rect 22112 27529 22140 27560
rect 22189 27557 22201 27591
rect 22235 27557 22247 27591
rect 22189 27551 22247 27557
rect 22097 27523 22155 27529
rect 22097 27489 22109 27523
rect 22143 27489 22155 27523
rect 22097 27483 22155 27489
rect 21637 27455 21695 27461
rect 21637 27452 21649 27455
rect 20916 27424 21649 27452
rect 21637 27421 21649 27424
rect 21683 27421 21695 27455
rect 21637 27415 21695 27421
rect 21818 27412 21824 27464
rect 21876 27412 21882 27464
rect 22370 27412 22376 27464
rect 22428 27412 22434 27464
rect 21174 27384 21180 27396
rect 20640 27356 21180 27384
rect 19582 27347 19640 27353
rect 21174 27344 21180 27356
rect 21232 27344 21238 27396
rect 21542 27344 21548 27396
rect 21600 27384 21606 27396
rect 22557 27387 22615 27393
rect 22557 27384 22569 27387
rect 21600 27356 22569 27384
rect 21600 27344 21606 27356
rect 22557 27353 22569 27356
rect 22603 27353 22615 27387
rect 22557 27347 22615 27353
rect 13633 27319 13691 27325
rect 13633 27285 13645 27319
rect 13679 27316 13691 27319
rect 13998 27316 14004 27328
rect 13679 27288 14004 27316
rect 13679 27285 13691 27288
rect 13633 27279 13691 27285
rect 13998 27276 14004 27288
rect 14056 27276 14062 27328
rect 17126 27276 17132 27328
rect 17184 27276 17190 27328
rect 19978 27276 19984 27328
rect 20036 27316 20042 27328
rect 20717 27319 20775 27325
rect 20717 27316 20729 27319
rect 20036 27288 20729 27316
rect 20036 27276 20042 27288
rect 20717 27285 20729 27288
rect 20763 27285 20775 27319
rect 20717 27279 20775 27285
rect 1104 27226 28888 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 28888 27226
rect 1104 27152 28888 27174
rect 12894 27072 12900 27124
rect 12952 27112 12958 27124
rect 13173 27115 13231 27121
rect 13173 27112 13185 27115
rect 12952 27084 13185 27112
rect 12952 27072 12958 27084
rect 13173 27081 13185 27084
rect 13219 27081 13231 27115
rect 13173 27075 13231 27081
rect 17678 27072 17684 27124
rect 17736 27072 17742 27124
rect 19058 27072 19064 27124
rect 19116 27072 19122 27124
rect 8938 27004 8944 27056
rect 8996 27044 9002 27056
rect 9186 27047 9244 27053
rect 9186 27044 9198 27047
rect 8996 27016 9198 27044
rect 8996 27004 9002 27016
rect 9186 27013 9198 27016
rect 9232 27013 9244 27047
rect 9186 27007 9244 27013
rect 12728 27016 14228 27044
rect 12728 26985 12756 27016
rect 14200 26988 14228 27016
rect 16942 27004 16948 27056
rect 17000 27044 17006 27056
rect 17494 27044 17500 27056
rect 17000 27016 17500 27044
rect 17000 27004 17006 27016
rect 17494 27004 17500 27016
rect 17552 27004 17558 27056
rect 20932 27047 20990 27053
rect 20932 27013 20944 27047
rect 20978 27044 20990 27047
rect 21542 27044 21548 27056
rect 20978 27016 21548 27044
rect 20978 27013 20990 27016
rect 20932 27007 20990 27013
rect 21542 27004 21548 27016
rect 21600 27004 21606 27056
rect 12713 26979 12771 26985
rect 12713 26945 12725 26979
rect 12759 26945 12771 26979
rect 12713 26939 12771 26945
rect 12986 26936 12992 26988
rect 13044 26976 13050 26988
rect 13541 26979 13599 26985
rect 13541 26976 13553 26979
rect 13044 26948 13553 26976
rect 13044 26936 13050 26948
rect 13541 26945 13553 26948
rect 13587 26945 13599 26979
rect 13541 26939 13599 26945
rect 13814 26936 13820 26988
rect 13872 26936 13878 26988
rect 13998 26936 14004 26988
rect 14056 26936 14062 26988
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 8938 26868 8944 26920
rect 8996 26868 9002 26920
rect 12618 26868 12624 26920
rect 12676 26868 12682 26920
rect 13357 26911 13415 26917
rect 13357 26908 13369 26911
rect 13096 26880 13369 26908
rect 13096 26784 13124 26880
rect 13357 26877 13369 26880
rect 13403 26877 13415 26911
rect 13357 26871 13415 26877
rect 13449 26911 13507 26917
rect 13449 26877 13461 26911
rect 13495 26877 13507 26911
rect 13449 26871 13507 26877
rect 13170 26800 13176 26852
rect 13228 26840 13234 26852
rect 13464 26840 13492 26871
rect 13630 26868 13636 26920
rect 13688 26868 13694 26920
rect 13722 26868 13728 26920
rect 13780 26908 13786 26920
rect 14108 26908 14136 26939
rect 14182 26936 14188 26988
rect 14240 26936 14246 26988
rect 16850 26936 16856 26988
rect 16908 26976 16914 26988
rect 17313 26979 17371 26985
rect 17313 26976 17325 26979
rect 16908 26948 17325 26976
rect 16908 26936 16914 26948
rect 17313 26945 17325 26948
rect 17359 26945 17371 26979
rect 17313 26939 17371 26945
rect 17954 26936 17960 26988
rect 18012 26976 18018 26988
rect 19242 26976 19248 26988
rect 18012 26948 19248 26976
rect 18012 26936 18018 26948
rect 19242 26936 19248 26948
rect 19300 26976 19306 26988
rect 19613 26979 19671 26985
rect 19613 26976 19625 26979
rect 19300 26948 19625 26976
rect 19300 26936 19306 26948
rect 19613 26945 19625 26948
rect 19659 26976 19671 26979
rect 19978 26976 19984 26988
rect 19659 26948 19984 26976
rect 19659 26945 19671 26948
rect 19613 26939 19671 26945
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 21174 26936 21180 26988
rect 21232 26936 21238 26988
rect 13780 26880 14136 26908
rect 13780 26868 13786 26880
rect 13228 26812 13492 26840
rect 13228 26800 13234 26812
rect 18230 26800 18236 26852
rect 18288 26840 18294 26852
rect 19797 26843 19855 26849
rect 19797 26840 19809 26843
rect 18288 26812 19809 26840
rect 18288 26800 18294 26812
rect 19797 26809 19809 26812
rect 19843 26809 19855 26843
rect 19797 26803 19855 26809
rect 10318 26732 10324 26784
rect 10376 26732 10382 26784
rect 13078 26732 13084 26784
rect 13136 26732 13142 26784
rect 14458 26732 14464 26784
rect 14516 26732 14522 26784
rect 19812 26772 19840 26803
rect 20806 26772 20812 26784
rect 19812 26744 20812 26772
rect 20806 26732 20812 26744
rect 20864 26732 20870 26784
rect 1104 26682 28888 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 28888 26682
rect 1104 26608 28888 26630
rect 13449 26571 13507 26577
rect 13449 26537 13461 26571
rect 13495 26568 13507 26571
rect 13630 26568 13636 26580
rect 13495 26540 13636 26568
rect 13495 26537 13507 26540
rect 13449 26531 13507 26537
rect 13630 26528 13636 26540
rect 13688 26528 13694 26580
rect 14182 26528 14188 26580
rect 14240 26568 14246 26580
rect 15749 26571 15807 26577
rect 15749 26568 15761 26571
rect 14240 26540 15761 26568
rect 14240 26528 14246 26540
rect 15749 26537 15761 26540
rect 15795 26537 15807 26571
rect 15749 26531 15807 26537
rect 13357 26503 13415 26509
rect 13357 26469 13369 26503
rect 13403 26500 13415 26503
rect 13817 26503 13875 26509
rect 13817 26500 13829 26503
rect 13403 26472 13829 26500
rect 13403 26469 13415 26472
rect 13357 26463 13415 26469
rect 13817 26469 13829 26472
rect 13863 26500 13875 26503
rect 13906 26500 13912 26512
rect 13863 26472 13912 26500
rect 13863 26469 13875 26472
rect 13817 26463 13875 26469
rect 13906 26460 13912 26472
rect 13964 26460 13970 26512
rect 15764 26500 15792 26531
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 19886 26568 19892 26580
rect 16724 26540 19892 26568
rect 16724 26528 16730 26540
rect 19886 26528 19892 26540
rect 19944 26528 19950 26580
rect 19978 26528 19984 26580
rect 20036 26528 20042 26580
rect 20441 26571 20499 26577
rect 20441 26537 20453 26571
rect 20487 26568 20499 26571
rect 21818 26568 21824 26580
rect 20487 26540 21824 26568
rect 20487 26537 20499 26540
rect 20441 26531 20499 26537
rect 21818 26528 21824 26540
rect 21876 26528 21882 26580
rect 17862 26500 17868 26512
rect 15764 26472 17868 26500
rect 17862 26460 17868 26472
rect 17920 26460 17926 26512
rect 19705 26503 19763 26509
rect 19705 26469 19717 26503
rect 19751 26500 19763 26503
rect 19794 26500 19800 26512
rect 19751 26472 19800 26500
rect 19751 26469 19763 26472
rect 19705 26463 19763 26469
rect 19794 26460 19800 26472
rect 19852 26460 19858 26512
rect 8938 26392 8944 26444
rect 8996 26432 9002 26444
rect 11977 26435 12035 26441
rect 11977 26432 11989 26435
rect 8996 26404 11989 26432
rect 8996 26392 9002 26404
rect 11977 26401 11989 26404
rect 12023 26401 12035 26435
rect 24486 26432 24492 26444
rect 11977 26395 12035 26401
rect 17972 26404 24492 26432
rect 12618 26324 12624 26376
rect 12676 26364 12682 26376
rect 13633 26367 13691 26373
rect 13633 26364 13645 26367
rect 12676 26336 13645 26364
rect 12676 26324 12682 26336
rect 13633 26333 13645 26336
rect 13679 26333 13691 26367
rect 13633 26327 13691 26333
rect 13909 26367 13967 26373
rect 13909 26333 13921 26367
rect 13955 26364 13967 26367
rect 14182 26364 14188 26376
rect 13955 26336 14188 26364
rect 13955 26333 13967 26336
rect 13909 26327 13967 26333
rect 14182 26324 14188 26336
rect 14240 26324 14246 26376
rect 14366 26324 14372 26376
rect 14424 26324 14430 26376
rect 14458 26324 14464 26376
rect 14516 26364 14522 26376
rect 17972 26373 18000 26404
rect 24486 26392 24492 26404
rect 24544 26392 24550 26444
rect 14625 26367 14683 26373
rect 14625 26364 14637 26367
rect 14516 26336 14637 26364
rect 14516 26324 14522 26336
rect 14625 26333 14637 26336
rect 14671 26333 14683 26367
rect 14625 26327 14683 26333
rect 17957 26367 18015 26373
rect 17957 26333 17969 26367
rect 18003 26333 18015 26367
rect 17957 26327 18015 26333
rect 19242 26324 19248 26376
rect 19300 26364 19306 26376
rect 19337 26367 19395 26373
rect 19337 26364 19349 26367
rect 19300 26336 19349 26364
rect 19300 26324 19306 26336
rect 19337 26333 19349 26336
rect 19383 26333 19395 26367
rect 19337 26327 19395 26333
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26364 19579 26367
rect 19567 26336 19932 26364
rect 19567 26333 19579 26336
rect 19521 26327 19579 26333
rect 12250 26305 12256 26308
rect 12244 26259 12256 26305
rect 12250 26256 12256 26259
rect 12308 26256 12314 26308
rect 18966 26256 18972 26308
rect 19024 26296 19030 26308
rect 19536 26296 19564 26327
rect 19024 26268 19564 26296
rect 19024 26256 19030 26268
rect 19610 26256 19616 26308
rect 19668 26296 19674 26308
rect 19797 26299 19855 26305
rect 19797 26296 19809 26299
rect 19668 26268 19809 26296
rect 19668 26256 19674 26268
rect 19797 26265 19809 26268
rect 19843 26265 19855 26299
rect 19904 26296 19932 26336
rect 20254 26324 20260 26376
rect 20312 26324 20318 26376
rect 20441 26367 20499 26373
rect 20441 26333 20453 26367
rect 20487 26364 20499 26367
rect 20898 26364 20904 26376
rect 20487 26336 20904 26364
rect 20487 26333 20499 26336
rect 20441 26327 20499 26333
rect 19997 26299 20055 26305
rect 19997 26296 20009 26299
rect 19904 26268 20009 26296
rect 19797 26259 19855 26265
rect 19997 26265 20009 26268
rect 20043 26265 20055 26299
rect 20456 26296 20484 26327
rect 20898 26324 20904 26336
rect 20956 26324 20962 26376
rect 19997 26259 20055 26265
rect 20180 26268 20484 26296
rect 12342 26188 12348 26240
rect 12400 26228 12406 26240
rect 12986 26228 12992 26240
rect 12400 26200 12992 26228
rect 12400 26188 12406 26200
rect 12986 26188 12992 26200
rect 13044 26188 13050 26240
rect 20180 26237 20208 26268
rect 20165 26231 20223 26237
rect 20165 26197 20177 26231
rect 20211 26197 20223 26231
rect 20165 26191 20223 26197
rect 1104 26138 28888 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 28888 26138
rect 1104 26064 28888 26086
rect 9217 26027 9275 26033
rect 9217 25993 9229 26027
rect 9263 26024 9275 26027
rect 9490 26024 9496 26036
rect 9263 25996 9496 26024
rect 9263 25993 9275 25996
rect 9217 25987 9275 25993
rect 9490 25984 9496 25996
rect 9548 25984 9554 26036
rect 12250 25984 12256 26036
rect 12308 25984 12314 26036
rect 13170 26024 13176 26036
rect 12406 25996 13176 26024
rect 12406 25900 12434 25996
rect 13170 25984 13176 25996
rect 13228 25984 13234 26036
rect 13446 25984 13452 26036
rect 13504 26024 13510 26036
rect 13541 26027 13599 26033
rect 13541 26024 13553 26027
rect 13504 25996 13553 26024
rect 13504 25984 13510 25996
rect 13541 25993 13553 25996
rect 13587 25993 13599 26027
rect 13541 25987 13599 25993
rect 16669 26027 16727 26033
rect 16669 25993 16681 26027
rect 16715 26024 16727 26027
rect 17586 26024 17592 26036
rect 16715 25996 17592 26024
rect 16715 25993 16727 25996
rect 16669 25987 16727 25993
rect 17586 25984 17592 25996
rect 17644 25984 17650 26036
rect 13909 25959 13967 25965
rect 13909 25956 13921 25959
rect 12728 25928 13921 25956
rect 9398 25848 9404 25900
rect 9456 25848 9462 25900
rect 9585 25891 9643 25897
rect 9585 25857 9597 25891
rect 9631 25888 9643 25891
rect 9858 25888 9864 25900
rect 9631 25860 9864 25888
rect 9631 25857 9643 25860
rect 9585 25851 9643 25857
rect 9858 25848 9864 25860
rect 9916 25888 9922 25900
rect 10318 25888 10324 25900
rect 9916 25860 10324 25888
rect 9916 25848 9922 25860
rect 10318 25848 10324 25860
rect 10376 25848 10382 25900
rect 11977 25891 12035 25897
rect 11977 25857 11989 25891
rect 12023 25888 12035 25891
rect 12406 25888 12440 25900
rect 12023 25860 12440 25888
rect 12023 25857 12035 25860
rect 11977 25851 12035 25857
rect 12434 25848 12440 25860
rect 12492 25848 12498 25900
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25857 12587 25891
rect 12529 25851 12587 25857
rect 11793 25823 11851 25829
rect 11793 25789 11805 25823
rect 11839 25820 11851 25823
rect 12250 25820 12256 25832
rect 11839 25792 12256 25820
rect 11839 25789 11851 25792
rect 11793 25783 11851 25789
rect 12250 25780 12256 25792
rect 12308 25780 12314 25832
rect 12342 25780 12348 25832
rect 12400 25820 12406 25832
rect 12544 25820 12572 25851
rect 12618 25848 12624 25900
rect 12676 25848 12682 25900
rect 12728 25897 12756 25928
rect 13909 25925 13921 25928
rect 13955 25925 13967 25959
rect 16758 25956 16764 25968
rect 13909 25919 13967 25925
rect 16224 25928 16764 25956
rect 12713 25891 12771 25897
rect 12713 25857 12725 25891
rect 12759 25857 12771 25891
rect 12713 25851 12771 25857
rect 12894 25848 12900 25900
rect 12952 25848 12958 25900
rect 12986 25848 12992 25900
rect 13044 25888 13050 25900
rect 13173 25891 13231 25897
rect 13173 25888 13185 25891
rect 13044 25860 13185 25888
rect 13044 25848 13050 25860
rect 13173 25857 13185 25860
rect 13219 25857 13231 25891
rect 13173 25851 13231 25857
rect 13633 25891 13691 25897
rect 13633 25857 13645 25891
rect 13679 25857 13691 25891
rect 13633 25851 13691 25857
rect 12400 25792 12572 25820
rect 12400 25780 12406 25792
rect 13078 25780 13084 25832
rect 13136 25780 13142 25832
rect 13648 25752 13676 25851
rect 16114 25848 16120 25900
rect 16172 25848 16178 25900
rect 16224 25897 16252 25928
rect 16758 25916 16764 25928
rect 16816 25916 16822 25968
rect 16942 25916 16948 25968
rect 17000 25916 17006 25968
rect 17037 25959 17095 25965
rect 17037 25925 17049 25959
rect 17083 25956 17095 25959
rect 17957 25959 18015 25965
rect 17957 25956 17969 25959
rect 17083 25928 17969 25956
rect 17083 25925 17095 25928
rect 17037 25919 17095 25925
rect 17957 25925 17969 25928
rect 18003 25925 18015 25959
rect 17957 25919 18015 25925
rect 16209 25891 16267 25897
rect 16209 25857 16221 25891
rect 16255 25857 16267 25891
rect 16209 25851 16267 25857
rect 16298 25848 16304 25900
rect 16356 25848 16362 25900
rect 16850 25897 16856 25900
rect 16848 25888 16856 25897
rect 16811 25860 16856 25888
rect 16848 25851 16856 25860
rect 16850 25848 16856 25851
rect 16908 25848 16914 25900
rect 17218 25848 17224 25900
rect 17276 25848 17282 25900
rect 17313 25891 17371 25897
rect 17313 25857 17325 25891
rect 17359 25857 17371 25891
rect 17313 25851 17371 25857
rect 13722 25780 13728 25832
rect 13780 25820 13786 25832
rect 13909 25823 13967 25829
rect 13909 25820 13921 25823
rect 13780 25792 13921 25820
rect 13780 25780 13786 25792
rect 13909 25789 13921 25792
rect 13955 25789 13967 25823
rect 17328 25820 17356 25851
rect 17862 25848 17868 25900
rect 17920 25888 17926 25900
rect 18171 25891 18229 25897
rect 18171 25888 18183 25891
rect 17920 25860 18183 25888
rect 17920 25848 17926 25860
rect 18171 25857 18183 25860
rect 18217 25857 18229 25891
rect 18171 25851 18229 25857
rect 18325 25891 18383 25897
rect 18325 25857 18337 25891
rect 18371 25857 18383 25891
rect 18325 25851 18383 25857
rect 17405 25823 17463 25829
rect 17405 25820 17417 25823
rect 17328 25792 17417 25820
rect 13909 25783 13967 25789
rect 17405 25789 17417 25792
rect 17451 25789 17463 25823
rect 17405 25783 17463 25789
rect 12176 25724 13676 25752
rect 17589 25755 17647 25761
rect 12176 25696 12204 25724
rect 17589 25721 17601 25755
rect 17635 25752 17647 25755
rect 18340 25752 18368 25851
rect 19426 25752 19432 25764
rect 17635 25724 19432 25752
rect 17635 25721 17647 25724
rect 17589 25715 17647 25721
rect 19426 25712 19432 25724
rect 19484 25712 19490 25764
rect 12158 25644 12164 25696
rect 12216 25644 12222 25696
rect 12618 25644 12624 25696
rect 12676 25684 12682 25696
rect 13630 25684 13636 25696
rect 12676 25656 13636 25684
rect 12676 25644 12682 25656
rect 13630 25644 13636 25656
rect 13688 25644 13694 25696
rect 13722 25644 13728 25696
rect 13780 25644 13786 25696
rect 15930 25644 15936 25696
rect 15988 25644 15994 25696
rect 1104 25594 28888 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 28888 25594
rect 1104 25520 28888 25542
rect 12437 25483 12495 25489
rect 12437 25449 12449 25483
rect 12483 25480 12495 25483
rect 13722 25480 13728 25492
rect 12483 25452 13728 25480
rect 12483 25449 12495 25452
rect 12437 25443 12495 25449
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 12986 25372 12992 25424
rect 13044 25372 13050 25424
rect 13170 25372 13176 25424
rect 13228 25412 13234 25424
rect 13265 25415 13323 25421
rect 13265 25412 13277 25415
rect 13228 25384 13277 25412
rect 13228 25372 13234 25384
rect 13265 25381 13277 25384
rect 13311 25412 13323 25415
rect 13630 25412 13636 25424
rect 13311 25384 13636 25412
rect 13311 25381 13323 25384
rect 13265 25375 13323 25381
rect 13630 25372 13636 25384
rect 13688 25372 13694 25424
rect 6825 25347 6883 25353
rect 6825 25313 6837 25347
rect 6871 25344 6883 25347
rect 8386 25344 8392 25356
rect 6871 25316 8392 25344
rect 6871 25313 6883 25316
rect 6825 25307 6883 25313
rect 8386 25304 8392 25316
rect 8444 25344 8450 25356
rect 8754 25344 8760 25356
rect 8444 25316 8760 25344
rect 8444 25304 8450 25316
rect 8754 25304 8760 25316
rect 8812 25304 8818 25356
rect 12158 25304 12164 25356
rect 12216 25344 12222 25356
rect 12216 25316 12848 25344
rect 12216 25304 12222 25316
rect 7006 25236 7012 25288
rect 7064 25236 7070 25288
rect 12250 25236 12256 25288
rect 12308 25236 12314 25288
rect 12434 25236 12440 25288
rect 12492 25236 12498 25288
rect 12526 25236 12532 25288
rect 12584 25236 12590 25288
rect 12820 25285 12848 25316
rect 12894 25304 12900 25356
rect 12952 25344 12958 25356
rect 13814 25344 13820 25356
rect 12952 25316 13820 25344
rect 12952 25304 12958 25316
rect 13814 25304 13820 25316
rect 13872 25304 13878 25356
rect 12805 25279 12863 25285
rect 12805 25245 12817 25279
rect 12851 25245 12863 25279
rect 12805 25239 12863 25245
rect 13081 25279 13139 25285
rect 13081 25245 13093 25279
rect 13127 25276 13139 25279
rect 13262 25276 13268 25288
rect 13127 25248 13268 25276
rect 13127 25245 13139 25248
rect 13081 25239 13139 25245
rect 13262 25236 13268 25248
rect 13320 25236 13326 25288
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 16025 25279 16083 25285
rect 16025 25276 16037 25279
rect 15436 25248 16037 25276
rect 15436 25236 15442 25248
rect 16025 25245 16037 25248
rect 16071 25276 16083 25279
rect 16114 25276 16120 25288
rect 16071 25248 16120 25276
rect 16071 25245 16083 25248
rect 16025 25239 16083 25245
rect 16114 25236 16120 25248
rect 16172 25236 16178 25288
rect 16209 25279 16267 25285
rect 16209 25245 16221 25279
rect 16255 25276 16267 25279
rect 17126 25276 17132 25288
rect 16255 25248 17132 25276
rect 16255 25245 16267 25248
rect 16209 25239 16267 25245
rect 17126 25236 17132 25248
rect 17184 25236 17190 25288
rect 6580 25211 6638 25217
rect 6580 25177 6592 25211
rect 6626 25208 6638 25211
rect 7834 25208 7840 25220
rect 6626 25180 7840 25208
rect 6626 25177 6638 25180
rect 6580 25171 6638 25177
rect 7834 25168 7840 25180
rect 7892 25168 7898 25220
rect 12621 25211 12679 25217
rect 12621 25177 12633 25211
rect 12667 25208 12679 25211
rect 13906 25208 13912 25220
rect 12667 25180 13912 25208
rect 12667 25177 12679 25180
rect 12621 25171 12679 25177
rect 5445 25143 5503 25149
rect 5445 25109 5457 25143
rect 5491 25140 5503 25143
rect 6362 25140 6368 25152
rect 5491 25112 6368 25140
rect 5491 25109 5503 25112
rect 5445 25103 5503 25109
rect 6362 25100 6368 25112
rect 6420 25100 6426 25152
rect 7561 25143 7619 25149
rect 7561 25109 7573 25143
rect 7607 25140 7619 25143
rect 8110 25140 8116 25152
rect 7607 25112 8116 25140
rect 7607 25109 7619 25112
rect 7561 25103 7619 25109
rect 8110 25100 8116 25112
rect 8168 25100 8174 25152
rect 12342 25100 12348 25152
rect 12400 25140 12406 25152
rect 12636 25140 12664 25171
rect 13906 25168 13912 25180
rect 13964 25168 13970 25220
rect 12400 25112 12664 25140
rect 12400 25100 12406 25112
rect 15654 25100 15660 25152
rect 15712 25140 15718 25152
rect 16117 25143 16175 25149
rect 16117 25140 16129 25143
rect 15712 25112 16129 25140
rect 15712 25100 15718 25112
rect 16117 25109 16129 25112
rect 16163 25109 16175 25143
rect 16117 25103 16175 25109
rect 1104 25050 28888 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 28888 25050
rect 1104 24976 28888 24998
rect 12526 24896 12532 24948
rect 12584 24936 12590 24948
rect 13538 24936 13544 24948
rect 12584 24908 13544 24936
rect 12584 24896 12590 24908
rect 13538 24896 13544 24908
rect 13596 24936 13602 24948
rect 13725 24939 13783 24945
rect 13725 24936 13737 24939
rect 13596 24908 13737 24936
rect 13596 24896 13602 24908
rect 13725 24905 13737 24908
rect 13771 24905 13783 24939
rect 13725 24899 13783 24905
rect 9024 24871 9082 24877
rect 3160 24840 3648 24868
rect 842 24760 848 24812
rect 900 24800 906 24812
rect 3160 24809 3188 24840
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 900 24772 1409 24800
rect 900 24760 906 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 2685 24803 2743 24809
rect 2685 24769 2697 24803
rect 2731 24769 2743 24803
rect 2685 24763 2743 24769
rect 3145 24803 3203 24809
rect 3145 24769 3157 24803
rect 3191 24769 3203 24803
rect 3412 24803 3470 24809
rect 3412 24798 3424 24803
rect 3145 24763 3203 24769
rect 3252 24770 3424 24798
rect 2498 24692 2504 24744
rect 2556 24692 2562 24744
rect 1581 24667 1639 24673
rect 1581 24633 1593 24667
rect 1627 24664 1639 24667
rect 2700 24664 2728 24763
rect 2869 24735 2927 24741
rect 2869 24701 2881 24735
rect 2915 24732 2927 24735
rect 3252 24732 3280 24770
rect 3412 24769 3424 24770
rect 3458 24769 3470 24803
rect 3620 24800 3648 24840
rect 9024 24837 9036 24871
rect 9070 24868 9082 24871
rect 9490 24868 9496 24880
rect 9070 24840 9496 24868
rect 9070 24837 9082 24840
rect 9024 24831 9082 24837
rect 9490 24828 9496 24840
rect 9548 24828 9554 24880
rect 16850 24828 16856 24880
rect 16908 24868 16914 24880
rect 19610 24868 19616 24880
rect 16908 24840 19616 24868
rect 16908 24828 16914 24840
rect 19610 24828 19616 24840
rect 19668 24828 19674 24880
rect 4706 24800 4712 24812
rect 3620 24772 4712 24800
rect 3412 24763 3470 24769
rect 4706 24760 4712 24772
rect 4764 24760 4770 24812
rect 4798 24760 4804 24812
rect 4856 24800 4862 24812
rect 4965 24803 5023 24809
rect 4965 24800 4977 24803
rect 4856 24772 4977 24800
rect 4856 24760 4862 24772
rect 4965 24769 4977 24772
rect 5011 24769 5023 24803
rect 4965 24763 5023 24769
rect 7466 24760 7472 24812
rect 7524 24809 7530 24812
rect 7524 24763 7536 24809
rect 7524 24760 7530 24763
rect 13354 24760 13360 24812
rect 13412 24800 13418 24812
rect 13541 24803 13599 24809
rect 13541 24800 13553 24803
rect 13412 24772 13553 24800
rect 13412 24760 13418 24772
rect 13541 24769 13553 24772
rect 13587 24769 13599 24803
rect 13541 24763 13599 24769
rect 13906 24760 13912 24812
rect 13964 24760 13970 24812
rect 2915 24704 3280 24732
rect 7745 24735 7803 24741
rect 2915 24701 2927 24704
rect 2869 24695 2927 24701
rect 7745 24701 7757 24735
rect 7791 24732 7803 24735
rect 8386 24732 8392 24744
rect 7791 24704 8392 24732
rect 7791 24701 7803 24704
rect 7745 24695 7803 24701
rect 8386 24692 8392 24704
rect 8444 24732 8450 24744
rect 8757 24735 8815 24741
rect 8757 24732 8769 24735
rect 8444 24704 8769 24732
rect 8444 24692 8450 24704
rect 8757 24701 8769 24704
rect 8803 24701 8815 24735
rect 8757 24695 8815 24701
rect 1627 24636 2728 24664
rect 1627 24633 1639 24636
rect 1581 24627 1639 24633
rect 13630 24624 13636 24676
rect 13688 24664 13694 24676
rect 14001 24667 14059 24673
rect 14001 24664 14013 24667
rect 13688 24636 14013 24664
rect 13688 24624 13694 24636
rect 14001 24633 14013 24636
rect 14047 24633 14059 24667
rect 14001 24627 14059 24633
rect 4525 24599 4583 24605
rect 4525 24565 4537 24599
rect 4571 24596 4583 24599
rect 5442 24596 5448 24608
rect 4571 24568 5448 24596
rect 4571 24565 4583 24568
rect 4525 24559 4583 24565
rect 5442 24556 5448 24568
rect 5500 24556 5506 24608
rect 6086 24556 6092 24608
rect 6144 24556 6150 24608
rect 6365 24599 6423 24605
rect 6365 24565 6377 24599
rect 6411 24596 6423 24599
rect 7006 24596 7012 24608
rect 6411 24568 7012 24596
rect 6411 24565 6423 24568
rect 6365 24559 6423 24565
rect 7006 24556 7012 24568
rect 7064 24556 7070 24608
rect 10134 24556 10140 24608
rect 10192 24556 10198 24608
rect 1104 24506 28888 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 28888 24506
rect 1104 24432 28888 24454
rect 4798 24352 4804 24404
rect 4856 24352 4862 24404
rect 5442 24352 5448 24404
rect 5500 24392 5506 24404
rect 6730 24392 6736 24404
rect 5500 24364 6736 24392
rect 5500 24352 5506 24364
rect 6730 24352 6736 24364
rect 6788 24392 6794 24404
rect 7285 24395 7343 24401
rect 7285 24392 7297 24395
rect 6788 24364 7297 24392
rect 6788 24352 6794 24364
rect 7285 24361 7297 24364
rect 7331 24361 7343 24395
rect 7285 24355 7343 24361
rect 7834 24352 7840 24404
rect 7892 24352 7898 24404
rect 6362 24284 6368 24336
rect 6420 24324 6426 24336
rect 6420 24296 7420 24324
rect 6420 24284 6426 24296
rect 4433 24259 4491 24265
rect 4433 24225 4445 24259
rect 4479 24256 4491 24259
rect 4893 24259 4951 24265
rect 4893 24256 4905 24259
rect 4479 24228 4905 24256
rect 4479 24225 4491 24228
rect 4433 24219 4491 24225
rect 4893 24225 4905 24228
rect 4939 24225 4951 24259
rect 4893 24219 4951 24225
rect 5442 24216 5448 24268
rect 5500 24216 5506 24268
rect 6086 24216 6092 24268
rect 6144 24256 6150 24268
rect 7392 24265 7420 24296
rect 12434 24284 12440 24336
rect 12492 24324 12498 24336
rect 13265 24327 13323 24333
rect 13265 24324 13277 24327
rect 12492 24296 13277 24324
rect 12492 24284 12498 24296
rect 13265 24293 13277 24296
rect 13311 24293 13323 24327
rect 13265 24287 13323 24293
rect 6549 24259 6607 24265
rect 6549 24256 6561 24259
rect 6144 24228 6561 24256
rect 6144 24216 6150 24228
rect 6549 24225 6561 24228
rect 6595 24256 6607 24259
rect 7377 24259 7435 24265
rect 6595 24228 6914 24256
rect 6595 24225 6607 24228
rect 6549 24219 6607 24225
rect 2498 24148 2504 24200
rect 2556 24188 2562 24200
rect 4617 24191 4675 24197
rect 4617 24188 4629 24191
rect 2556 24160 4629 24188
rect 2556 24148 2562 24160
rect 4617 24157 4629 24160
rect 4663 24188 4675 24191
rect 5902 24188 5908 24200
rect 4663 24160 5908 24188
rect 4663 24157 4675 24160
rect 4617 24151 4675 24157
rect 5902 24148 5908 24160
rect 5960 24148 5966 24200
rect 6362 24148 6368 24200
rect 6420 24148 6426 24200
rect 6886 24188 6914 24228
rect 7377 24225 7389 24259
rect 7423 24225 7435 24259
rect 8294 24256 8300 24268
rect 7377 24219 7435 24225
rect 8036 24228 8300 24256
rect 8036 24197 8064 24228
rect 8294 24216 8300 24228
rect 8352 24256 8358 24268
rect 9398 24256 9404 24268
rect 8352 24228 9404 24256
rect 8352 24216 8358 24228
rect 9398 24216 9404 24228
rect 9456 24216 9462 24268
rect 13538 24216 13544 24268
rect 13596 24216 13602 24268
rect 7561 24191 7619 24197
rect 7561 24188 7573 24191
rect 6886 24160 7573 24188
rect 7561 24157 7573 24160
rect 7607 24157 7619 24191
rect 7561 24151 7619 24157
rect 8021 24191 8079 24197
rect 8021 24157 8033 24191
rect 8067 24157 8079 24191
rect 8021 24151 8079 24157
rect 8110 24148 8116 24200
rect 8168 24148 8174 24200
rect 13630 24148 13636 24200
rect 13688 24148 13694 24200
rect 7006 24080 7012 24132
rect 7064 24120 7070 24132
rect 7282 24120 7288 24132
rect 7064 24092 7288 24120
rect 7064 24080 7070 24092
rect 7282 24080 7288 24092
rect 7340 24080 7346 24132
rect 5813 24055 5871 24061
rect 5813 24021 5825 24055
rect 5859 24052 5871 24055
rect 5994 24052 6000 24064
rect 5859 24024 6000 24052
rect 5859 24021 5871 24024
rect 5813 24015 5871 24021
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 7190 24012 7196 24064
rect 7248 24012 7254 24064
rect 7742 24012 7748 24064
rect 7800 24012 7806 24064
rect 1104 23962 28888 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 28888 23962
rect 1104 23888 28888 23910
rect 6362 23808 6368 23860
rect 6420 23848 6426 23860
rect 6549 23851 6607 23857
rect 6549 23848 6561 23851
rect 6420 23820 6561 23848
rect 6420 23808 6426 23820
rect 6549 23817 6561 23820
rect 6595 23817 6607 23851
rect 7466 23848 7472 23860
rect 6549 23811 6607 23817
rect 6886 23820 7472 23848
rect 6457 23783 6515 23789
rect 6457 23749 6469 23783
rect 6503 23780 6515 23783
rect 6886 23780 6914 23820
rect 7466 23808 7472 23820
rect 7524 23808 7530 23860
rect 16301 23851 16359 23857
rect 15304 23820 16068 23848
rect 6503 23752 6914 23780
rect 6503 23749 6515 23752
rect 6457 23743 6515 23749
rect 10134 23740 10140 23792
rect 10192 23780 10198 23792
rect 10229 23783 10287 23789
rect 10229 23780 10241 23783
rect 10192 23752 10241 23780
rect 10192 23740 10198 23752
rect 10229 23749 10241 23752
rect 10275 23749 10287 23783
rect 10229 23743 10287 23749
rect 15304 23724 15332 23820
rect 15396 23752 15884 23780
rect 5902 23672 5908 23724
rect 5960 23672 5966 23724
rect 5994 23672 6000 23724
rect 6052 23672 6058 23724
rect 6730 23672 6736 23724
rect 6788 23672 6794 23724
rect 7190 23672 7196 23724
rect 7248 23672 7254 23724
rect 7285 23715 7343 23721
rect 7285 23681 7297 23715
rect 7331 23712 7343 23715
rect 8294 23712 8300 23724
rect 7331 23684 8300 23712
rect 7331 23681 7343 23684
rect 7285 23675 7343 23681
rect 5920 23576 5948 23672
rect 6362 23604 6368 23656
rect 6420 23604 6426 23656
rect 6822 23604 6828 23656
rect 6880 23604 6886 23656
rect 7300 23576 7328 23675
rect 8294 23672 8300 23684
rect 8352 23672 8358 23724
rect 9766 23672 9772 23724
rect 9824 23672 9830 23724
rect 10410 23672 10416 23724
rect 10468 23672 10474 23724
rect 13630 23672 13636 23724
rect 13688 23712 13694 23724
rect 15013 23715 15071 23721
rect 15013 23712 15025 23715
rect 13688 23684 15025 23712
rect 13688 23672 13694 23684
rect 15013 23681 15025 23684
rect 15059 23681 15071 23715
rect 15013 23675 15071 23681
rect 9858 23604 9864 23656
rect 9916 23604 9922 23656
rect 5920 23548 7328 23576
rect 10137 23579 10195 23585
rect 10137 23545 10149 23579
rect 10183 23576 10195 23579
rect 11422 23576 11428 23588
rect 10183 23548 11428 23576
rect 10183 23545 10195 23548
rect 10137 23539 10195 23545
rect 11422 23536 11428 23548
rect 11480 23536 11486 23588
rect 15028 23576 15056 23675
rect 15286 23672 15292 23724
rect 15344 23672 15350 23724
rect 15396 23721 15424 23752
rect 15381 23715 15439 23721
rect 15381 23681 15393 23715
rect 15427 23681 15439 23715
rect 15381 23675 15439 23681
rect 15654 23672 15660 23724
rect 15712 23672 15718 23724
rect 15746 23672 15752 23724
rect 15804 23672 15810 23724
rect 15856 23712 15884 23752
rect 15930 23740 15936 23792
rect 15988 23740 15994 23792
rect 16040 23789 16068 23820
rect 16301 23817 16313 23851
rect 16347 23848 16359 23851
rect 16347 23820 16896 23848
rect 16347 23817 16359 23820
rect 16301 23811 16359 23817
rect 16868 23789 16896 23820
rect 17218 23808 17224 23860
rect 17276 23808 17282 23860
rect 18966 23808 18972 23860
rect 19024 23848 19030 23860
rect 19245 23851 19303 23857
rect 19245 23848 19257 23851
rect 19024 23820 19257 23848
rect 19024 23808 19030 23820
rect 19245 23817 19257 23820
rect 19291 23848 19303 23851
rect 19291 23820 19748 23848
rect 19291 23817 19303 23820
rect 19245 23811 19303 23817
rect 16025 23783 16083 23789
rect 16025 23749 16037 23783
rect 16071 23749 16083 23783
rect 16025 23743 16083 23749
rect 16853 23783 16911 23789
rect 16853 23749 16865 23783
rect 16899 23749 16911 23783
rect 16853 23743 16911 23749
rect 18138 23740 18144 23792
rect 18196 23780 18202 23792
rect 19397 23783 19455 23789
rect 19397 23780 19409 23783
rect 18196 23752 19409 23780
rect 18196 23740 18202 23752
rect 19397 23749 19409 23752
rect 19443 23749 19455 23783
rect 19397 23743 19455 23749
rect 19610 23740 19616 23792
rect 19668 23740 19674 23792
rect 16114 23712 16120 23724
rect 16172 23721 16178 23724
rect 19720 23721 19748 23820
rect 15856 23684 16120 23712
rect 16114 23672 16120 23684
rect 16172 23675 16180 23721
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 16945 23715 17003 23721
rect 16945 23681 16957 23715
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23681 17095 23715
rect 17037 23675 17095 23681
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23681 19763 23715
rect 19705 23675 19763 23681
rect 19889 23715 19947 23721
rect 19889 23681 19901 23715
rect 19935 23681 19947 23715
rect 19889 23675 19947 23681
rect 16172 23672 16178 23675
rect 15565 23647 15623 23653
rect 15565 23613 15577 23647
rect 15611 23644 15623 23647
rect 16684 23644 16712 23675
rect 15611 23616 16712 23644
rect 15611 23613 15623 23616
rect 15565 23607 15623 23613
rect 16960 23576 16988 23675
rect 15028 23548 16988 23576
rect 5718 23468 5724 23520
rect 5776 23468 5782 23520
rect 7009 23511 7067 23517
rect 7009 23477 7021 23511
rect 7055 23508 7067 23511
rect 7098 23508 7104 23520
rect 7055 23480 7104 23508
rect 7055 23477 7067 23480
rect 7009 23471 7067 23477
rect 7098 23468 7104 23480
rect 7156 23468 7162 23520
rect 10597 23511 10655 23517
rect 10597 23477 10609 23511
rect 10643 23508 10655 23511
rect 11238 23508 11244 23520
rect 10643 23480 11244 23508
rect 10643 23477 10655 23480
rect 10597 23471 10655 23477
rect 11238 23468 11244 23480
rect 11296 23468 11302 23520
rect 15105 23511 15163 23517
rect 15105 23477 15117 23511
rect 15151 23508 15163 23511
rect 16850 23508 16856 23520
rect 15151 23480 16856 23508
rect 15151 23477 15163 23480
rect 15105 23471 15163 23477
rect 16850 23468 16856 23480
rect 16908 23508 16914 23520
rect 17052 23508 17080 23675
rect 17954 23604 17960 23656
rect 18012 23644 18018 23656
rect 18966 23644 18972 23656
rect 18012 23616 18972 23644
rect 18012 23604 18018 23616
rect 18966 23604 18972 23616
rect 19024 23644 19030 23656
rect 19904 23644 19932 23675
rect 28258 23672 28264 23724
rect 28316 23672 28322 23724
rect 19024 23616 19932 23644
rect 19024 23604 19030 23616
rect 16908 23480 17080 23508
rect 16908 23468 16914 23480
rect 19426 23468 19432 23520
rect 19484 23468 19490 23520
rect 19702 23468 19708 23520
rect 19760 23468 19766 23520
rect 28442 23468 28448 23520
rect 28500 23468 28506 23520
rect 1104 23418 28888 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 28888 23418
rect 1104 23344 28888 23366
rect 10321 23307 10379 23313
rect 10321 23273 10333 23307
rect 10367 23304 10379 23307
rect 10410 23304 10416 23316
rect 10367 23276 10416 23304
rect 10367 23273 10379 23276
rect 10321 23267 10379 23273
rect 10410 23264 10416 23276
rect 10468 23304 10474 23316
rect 11425 23307 11483 23313
rect 10468 23276 10824 23304
rect 10468 23264 10474 23276
rect 4706 23128 4712 23180
rect 4764 23168 4770 23180
rect 5261 23171 5319 23177
rect 5261 23168 5273 23171
rect 4764 23140 5273 23168
rect 4764 23128 4770 23140
rect 5261 23137 5273 23140
rect 5307 23137 5319 23171
rect 5261 23131 5319 23137
rect 6288 23140 7420 23168
rect 5276 23100 5304 23131
rect 5350 23100 5356 23112
rect 5276 23072 5356 23100
rect 5350 23060 5356 23072
rect 5408 23100 5414 23112
rect 6288 23100 6316 23140
rect 5408 23072 6316 23100
rect 6733 23103 6791 23109
rect 5408 23060 5414 23072
rect 6733 23069 6745 23103
rect 6779 23100 6791 23103
rect 6822 23100 6828 23112
rect 6779 23072 6828 23100
rect 6779 23069 6791 23072
rect 6733 23063 6791 23069
rect 6822 23060 6828 23072
rect 6880 23060 6886 23112
rect 7098 23060 7104 23112
rect 7156 23060 7162 23112
rect 7392 23109 7420 23140
rect 9950 23128 9956 23180
rect 10008 23168 10014 23180
rect 10796 23177 10824 23276
rect 11425 23273 11437 23307
rect 11471 23304 11483 23307
rect 13262 23304 13268 23316
rect 11471 23276 13268 23304
rect 11471 23273 11483 23276
rect 11425 23267 11483 23273
rect 13262 23264 13268 23276
rect 13320 23264 13326 23316
rect 16850 23264 16856 23316
rect 16908 23264 16914 23316
rect 27709 23307 27767 23313
rect 27709 23273 27721 23307
rect 27755 23304 27767 23307
rect 28258 23304 28264 23316
rect 27755 23276 28264 23304
rect 27755 23273 27767 23276
rect 27709 23267 27767 23273
rect 28258 23264 28264 23276
rect 28316 23264 28322 23316
rect 12069 23239 12127 23245
rect 12069 23205 12081 23239
rect 12115 23236 12127 23239
rect 13354 23236 13360 23248
rect 12115 23208 13360 23236
rect 12115 23205 12127 23208
rect 12069 23199 12127 23205
rect 13354 23196 13360 23208
rect 13412 23196 13418 23248
rect 17037 23239 17095 23245
rect 17037 23205 17049 23239
rect 17083 23236 17095 23239
rect 18138 23236 18144 23248
rect 17083 23208 18144 23236
rect 17083 23205 17095 23208
rect 17037 23199 17095 23205
rect 10689 23171 10747 23177
rect 10689 23168 10701 23171
rect 10008 23140 10701 23168
rect 10008 23128 10014 23140
rect 10689 23137 10701 23140
rect 10735 23137 10747 23171
rect 10689 23131 10747 23137
rect 10781 23171 10839 23177
rect 10781 23137 10793 23171
rect 10827 23137 10839 23171
rect 10781 23131 10839 23137
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23100 7435 23103
rect 8386 23100 8392 23112
rect 7423 23072 8392 23100
rect 7423 23069 7435 23072
rect 7377 23063 7435 23069
rect 8386 23060 8392 23072
rect 8444 23100 8450 23112
rect 8938 23100 8944 23112
rect 8444 23072 8944 23100
rect 8444 23060 8450 23072
rect 8938 23060 8944 23072
rect 8996 23060 9002 23112
rect 9766 23060 9772 23112
rect 9824 23100 9830 23112
rect 10413 23103 10471 23109
rect 10413 23100 10425 23103
rect 9824 23072 10425 23100
rect 9824 23060 9830 23072
rect 10413 23069 10425 23072
rect 10459 23069 10471 23103
rect 10413 23063 10471 23069
rect 10594 23060 10600 23112
rect 10652 23100 10658 23112
rect 11149 23103 11207 23109
rect 11149 23100 11161 23103
rect 10652 23072 11161 23100
rect 10652 23060 10658 23072
rect 11149 23069 11161 23072
rect 11195 23069 11207 23103
rect 11149 23063 11207 23069
rect 11238 23060 11244 23112
rect 11296 23060 11302 23112
rect 11422 23060 11428 23112
rect 11480 23060 11486 23112
rect 17144 23109 17172 23208
rect 18138 23196 18144 23208
rect 18196 23196 18202 23248
rect 19610 23196 19616 23248
rect 19668 23236 19674 23248
rect 19668 23208 20576 23236
rect 19668 23196 19674 23208
rect 17405 23171 17463 23177
rect 17405 23137 17417 23171
rect 17451 23168 17463 23171
rect 17954 23168 17960 23180
rect 17451 23140 17960 23168
rect 17451 23137 17463 23140
rect 17405 23131 17463 23137
rect 17954 23128 17960 23140
rect 18012 23128 18018 23180
rect 20548 23177 20576 23208
rect 18969 23171 19027 23177
rect 18969 23137 18981 23171
rect 19015 23168 19027 23171
rect 19981 23171 20039 23177
rect 19981 23168 19993 23171
rect 19015 23140 19993 23168
rect 19015 23137 19027 23140
rect 18969 23131 19027 23137
rect 19981 23137 19993 23140
rect 20027 23137 20039 23171
rect 19981 23131 20039 23137
rect 20533 23171 20591 23177
rect 20533 23137 20545 23171
rect 20579 23137 20591 23171
rect 20533 23131 20591 23137
rect 12161 23103 12219 23109
rect 12161 23100 12173 23103
rect 11716 23072 12173 23100
rect 11716 23044 11744 23072
rect 12161 23069 12173 23072
rect 12207 23069 12219 23103
rect 12161 23063 12219 23069
rect 17129 23103 17187 23109
rect 17129 23069 17141 23103
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 17221 23103 17279 23109
rect 17221 23069 17233 23103
rect 17267 23069 17279 23103
rect 17221 23063 17279 23069
rect 18693 23103 18751 23109
rect 18693 23069 18705 23103
rect 18739 23069 18751 23103
rect 18693 23063 18751 23069
rect 5528 23035 5586 23041
rect 5528 23001 5540 23035
rect 5574 23032 5586 23035
rect 5718 23032 5724 23044
rect 5574 23004 5724 23032
rect 5574 23001 5586 23004
rect 5528 22995 5586 23001
rect 5718 22992 5724 23004
rect 5776 22992 5782 23044
rect 6917 23035 6975 23041
rect 6917 23001 6929 23035
rect 6963 23001 6975 23035
rect 6917 22995 6975 23001
rect 6641 22967 6699 22973
rect 6641 22933 6653 22967
rect 6687 22964 6699 22967
rect 6730 22964 6736 22976
rect 6687 22936 6736 22964
rect 6687 22933 6699 22936
rect 6641 22927 6699 22933
rect 6730 22924 6736 22936
rect 6788 22924 6794 22976
rect 6932 22964 6960 22995
rect 7006 22992 7012 23044
rect 7064 22992 7070 23044
rect 7644 23035 7702 23041
rect 7644 23001 7656 23035
rect 7690 23032 7702 23035
rect 8110 23032 8116 23044
rect 7690 23004 8116 23032
rect 7690 23001 7702 23004
rect 7644 22995 7702 23001
rect 8110 22992 8116 23004
rect 8168 22992 8174 23044
rect 8662 22992 8668 23044
rect 8720 23032 8726 23044
rect 9186 23035 9244 23041
rect 9186 23032 9198 23035
rect 8720 23004 9198 23032
rect 8720 22992 8726 23004
rect 9186 23001 9198 23004
rect 9232 23001 9244 23035
rect 9186 22995 9244 23001
rect 10134 22992 10140 23044
rect 10192 23032 10198 23044
rect 10898 23035 10956 23041
rect 10898 23032 10910 23035
rect 10192 23004 10910 23032
rect 10192 22992 10198 23004
rect 10898 23001 10910 23004
rect 10944 23001 10956 23035
rect 10898 22995 10956 23001
rect 11698 22992 11704 23044
rect 11756 22992 11762 23044
rect 11885 23035 11943 23041
rect 11885 23001 11897 23035
rect 11931 23001 11943 23035
rect 11885 22995 11943 23001
rect 7098 22964 7104 22976
rect 6932 22936 7104 22964
rect 7098 22924 7104 22936
rect 7156 22924 7162 22976
rect 7285 22967 7343 22973
rect 7285 22933 7297 22967
rect 7331 22964 7343 22967
rect 7466 22964 7472 22976
rect 7331 22936 7472 22964
rect 7331 22933 7343 22936
rect 7285 22927 7343 22933
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 8754 22924 8760 22976
rect 8812 22924 8818 22976
rect 11057 22967 11115 22973
rect 11057 22933 11069 22967
rect 11103 22964 11115 22967
rect 11790 22964 11796 22976
rect 11103 22936 11796 22964
rect 11103 22933 11115 22936
rect 11057 22927 11115 22933
rect 11790 22924 11796 22936
rect 11848 22964 11854 22976
rect 11900 22964 11928 22995
rect 15746 22992 15752 23044
rect 15804 23032 15810 23044
rect 16669 23035 16727 23041
rect 16669 23032 16681 23035
rect 15804 23004 16681 23032
rect 15804 22992 15810 23004
rect 16669 23001 16681 23004
rect 16715 23001 16727 23035
rect 16669 22995 16727 23001
rect 16758 22992 16764 23044
rect 16816 23032 16822 23044
rect 17236 23032 17264 23063
rect 16816 23004 17264 23032
rect 18708 23032 18736 23063
rect 18874 23060 18880 23112
rect 18932 23060 18938 23112
rect 19426 23060 19432 23112
rect 19484 23100 19490 23112
rect 19797 23103 19855 23109
rect 19797 23100 19809 23103
rect 19484 23072 19809 23100
rect 19484 23060 19490 23072
rect 19797 23069 19809 23072
rect 19843 23069 19855 23103
rect 19797 23063 19855 23069
rect 27522 23060 27528 23112
rect 27580 23060 27586 23112
rect 19702 23032 19708 23044
rect 18708 23004 19708 23032
rect 16816 22992 16822 23004
rect 19702 22992 19708 23004
rect 19760 22992 19766 23044
rect 11848 22936 11928 22964
rect 11848 22924 11854 22936
rect 12342 22924 12348 22976
rect 12400 22924 12406 22976
rect 16114 22924 16120 22976
rect 16172 22964 16178 22976
rect 16869 22967 16927 22973
rect 16869 22964 16881 22967
rect 16172 22936 16881 22964
rect 16172 22924 16178 22936
rect 16869 22933 16881 22936
rect 16915 22933 16927 22967
rect 16869 22927 16927 22933
rect 17126 22924 17132 22976
rect 17184 22924 17190 22976
rect 18506 22924 18512 22976
rect 18564 22924 18570 22976
rect 19242 22924 19248 22976
rect 19300 22924 19306 22976
rect 1104 22874 28888 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 28888 22874
rect 1104 22800 28888 22822
rect 6362 22720 6368 22772
rect 6420 22720 6426 22772
rect 6730 22720 6736 22772
rect 6788 22760 6794 22772
rect 6914 22760 6920 22772
rect 6788 22732 6920 22760
rect 6788 22720 6794 22732
rect 6914 22720 6920 22732
rect 6972 22720 6978 22772
rect 8110 22720 8116 22772
rect 8168 22720 8174 22772
rect 10594 22720 10600 22772
rect 10652 22720 10658 22772
rect 14737 22763 14795 22769
rect 14737 22729 14749 22763
rect 14783 22760 14795 22763
rect 15286 22760 15292 22772
rect 14783 22732 15292 22760
rect 14783 22729 14795 22732
rect 14737 22723 14795 22729
rect 15286 22720 15292 22732
rect 15344 22720 15350 22772
rect 15746 22720 15752 22772
rect 15804 22760 15810 22772
rect 16022 22760 16028 22772
rect 15804 22732 16028 22760
rect 15804 22720 15810 22732
rect 16022 22720 16028 22732
rect 16080 22760 16086 22772
rect 16209 22763 16267 22769
rect 16209 22760 16221 22763
rect 16080 22732 16221 22760
rect 16080 22720 16086 22732
rect 16209 22729 16221 22732
rect 16255 22729 16267 22763
rect 19242 22760 19248 22772
rect 16209 22723 16267 22729
rect 17696 22732 19248 22760
rect 6549 22695 6607 22701
rect 6549 22661 6561 22695
rect 6595 22692 6607 22695
rect 6595 22664 6776 22692
rect 6595 22661 6607 22664
rect 6549 22655 6607 22661
rect 6748 22636 6776 22664
rect 6822 22652 6828 22704
rect 6880 22692 6886 22704
rect 8662 22692 8668 22704
rect 6880 22664 8668 22692
rect 6880 22652 6886 22664
rect 8662 22652 8668 22664
rect 8720 22652 8726 22704
rect 8754 22652 8760 22704
rect 8812 22692 8818 22704
rect 8812 22664 8984 22692
rect 8812 22652 8818 22664
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22593 6699 22627
rect 6641 22587 6699 22593
rect 6656 22556 6684 22587
rect 6730 22584 6736 22636
rect 6788 22584 6794 22636
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22624 6975 22627
rect 7282 22624 7288 22636
rect 6963 22596 7288 22624
rect 6963 22593 6975 22596
rect 6917 22587 6975 22593
rect 7282 22584 7288 22596
rect 7340 22584 7346 22636
rect 7466 22584 7472 22636
rect 7524 22584 7530 22636
rect 8294 22584 8300 22636
rect 8352 22624 8358 22636
rect 8956 22633 8984 22664
rect 10060 22664 10548 22692
rect 8849 22627 8907 22633
rect 8849 22624 8861 22627
rect 8352 22596 8861 22624
rect 8352 22584 8358 22596
rect 8849 22593 8861 22596
rect 8895 22593 8907 22627
rect 8849 22587 8907 22593
rect 8941 22627 8999 22633
rect 8941 22593 8953 22627
rect 8987 22624 8999 22627
rect 9766 22624 9772 22636
rect 8987 22596 9772 22624
rect 8987 22593 8999 22596
rect 8941 22587 8999 22593
rect 9766 22584 9772 22596
rect 9824 22624 9830 22636
rect 9861 22627 9919 22633
rect 9861 22624 9873 22627
rect 9824 22596 9873 22624
rect 9824 22584 9830 22596
rect 9861 22593 9873 22596
rect 9907 22593 9919 22627
rect 9861 22587 9919 22593
rect 9950 22584 9956 22636
rect 10008 22584 10014 22636
rect 10060 22633 10088 22664
rect 10520 22636 10548 22664
rect 10045 22627 10103 22633
rect 10045 22593 10057 22627
rect 10091 22593 10103 22627
rect 10045 22587 10103 22593
rect 10134 22584 10140 22636
rect 10192 22624 10198 22636
rect 10413 22627 10471 22633
rect 10413 22624 10425 22627
rect 10192 22596 10425 22624
rect 10192 22584 10198 22596
rect 10413 22593 10425 22596
rect 10459 22593 10471 22627
rect 10413 22587 10471 22593
rect 10502 22584 10508 22636
rect 10560 22624 10566 22636
rect 10597 22627 10655 22633
rect 10597 22624 10609 22627
rect 10560 22596 10609 22624
rect 10560 22584 10566 22596
rect 10597 22593 10609 22596
rect 10643 22593 10655 22627
rect 10597 22587 10655 22593
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 16114 22584 16120 22636
rect 16172 22584 16178 22636
rect 16393 22627 16451 22633
rect 16393 22593 16405 22627
rect 16439 22624 16451 22627
rect 16669 22627 16727 22633
rect 16669 22624 16681 22627
rect 16439 22596 16681 22624
rect 16439 22593 16451 22596
rect 16393 22587 16451 22593
rect 16669 22593 16681 22596
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 16850 22584 16856 22636
rect 16908 22624 16914 22636
rect 17696 22633 17724 22732
rect 19242 22720 19248 22732
rect 19300 22720 19306 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 19705 22763 19763 22769
rect 19705 22760 19717 22763
rect 19484 22732 19717 22760
rect 19484 22720 19490 22732
rect 19705 22729 19717 22732
rect 19751 22729 19763 22763
rect 19705 22723 19763 22729
rect 18248 22664 21128 22692
rect 17221 22627 17279 22633
rect 17221 22624 17233 22627
rect 16908 22596 17233 22624
rect 16908 22584 16914 22596
rect 17221 22593 17233 22596
rect 17267 22593 17279 22627
rect 17221 22587 17279 22593
rect 17681 22627 17739 22633
rect 17681 22593 17693 22627
rect 17727 22593 17739 22627
rect 17681 22587 17739 22593
rect 17954 22584 17960 22636
rect 18012 22584 18018 22636
rect 18046 22584 18052 22636
rect 18104 22624 18110 22636
rect 18248 22633 18276 22664
rect 18506 22633 18512 22636
rect 18233 22627 18291 22633
rect 18233 22624 18245 22627
rect 18104 22596 18245 22624
rect 18104 22584 18110 22596
rect 18233 22593 18245 22596
rect 18279 22593 18291 22627
rect 18500 22624 18512 22633
rect 18467 22596 18512 22624
rect 18233 22587 18291 22593
rect 18500 22587 18512 22596
rect 18506 22584 18512 22587
rect 18564 22584 18570 22636
rect 21100 22633 21128 22664
rect 20818 22627 20876 22633
rect 20818 22624 20830 22627
rect 19536 22596 20830 22624
rect 6822 22556 6828 22568
rect 6656 22528 6828 22556
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 10321 22559 10379 22565
rect 10321 22525 10333 22559
rect 10367 22556 10379 22559
rect 11698 22556 11704 22568
rect 10367 22528 11704 22556
rect 10367 22525 10379 22528
rect 10321 22519 10379 22525
rect 11698 22516 11704 22528
rect 11756 22516 11762 22568
rect 16574 22516 16580 22568
rect 16632 22556 16638 22568
rect 16868 22556 16896 22584
rect 16632 22528 16896 22556
rect 17773 22559 17831 22565
rect 16632 22516 16638 22528
rect 17773 22525 17785 22559
rect 17819 22556 17831 22559
rect 18138 22556 18144 22568
rect 17819 22528 18144 22556
rect 17819 22525 17831 22528
rect 17773 22519 17831 22525
rect 18138 22516 18144 22528
rect 18196 22516 18202 22568
rect 16393 22491 16451 22497
rect 16393 22457 16405 22491
rect 16439 22488 16451 22491
rect 16758 22488 16764 22500
rect 16439 22460 16764 22488
rect 16439 22457 16451 22460
rect 16393 22451 16451 22457
rect 16758 22448 16764 22460
rect 16816 22448 16822 22500
rect 18141 22423 18199 22429
rect 18141 22389 18153 22423
rect 18187 22420 18199 22423
rect 19536 22420 19564 22596
rect 20818 22593 20830 22596
rect 20864 22593 20876 22627
rect 20818 22587 20876 22593
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 28534 22516 28540 22568
rect 28592 22516 28598 22568
rect 19610 22448 19616 22500
rect 19668 22448 19674 22500
rect 18187 22392 19564 22420
rect 18187 22389 18199 22392
rect 18141 22383 18199 22389
rect 1104 22330 28888 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 28888 22330
rect 1104 22256 28888 22278
rect 7285 22219 7343 22225
rect 7285 22216 7297 22219
rect 6886 22188 7297 22216
rect 6886 22160 6914 22188
rect 7285 22185 7297 22188
rect 7331 22185 7343 22219
rect 7285 22179 7343 22185
rect 11793 22219 11851 22225
rect 11793 22185 11805 22219
rect 11839 22216 11851 22219
rect 12342 22216 12348 22228
rect 11839 22188 12348 22216
rect 11839 22185 11851 22188
rect 11793 22179 11851 22185
rect 12342 22176 12348 22188
rect 12400 22176 12406 22228
rect 12805 22219 12863 22225
rect 12805 22185 12817 22219
rect 12851 22185 12863 22219
rect 12805 22179 12863 22185
rect 6822 22108 6828 22160
rect 6880 22120 6914 22160
rect 6880 22108 6886 22120
rect 7098 22108 7104 22160
rect 7156 22108 7162 22160
rect 12820 22148 12848 22179
rect 18138 22176 18144 22228
rect 18196 22216 18202 22228
rect 18598 22216 18604 22228
rect 18196 22188 18604 22216
rect 18196 22176 18202 22188
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 18693 22219 18751 22225
rect 18693 22185 18705 22219
rect 18739 22216 18751 22219
rect 18874 22216 18880 22228
rect 18739 22188 18880 22216
rect 18739 22185 18751 22188
rect 18693 22179 18751 22185
rect 18874 22176 18880 22188
rect 18932 22176 18938 22228
rect 12452 22120 12848 22148
rect 6914 22040 6920 22092
rect 6972 22080 6978 22092
rect 11701 22083 11759 22089
rect 6972 22052 7328 22080
rect 6972 22040 6978 22052
rect 7300 22021 7328 22052
rect 11701 22049 11713 22083
rect 11747 22080 11759 22083
rect 11790 22080 11796 22092
rect 11747 22052 11796 22080
rect 11747 22049 11759 22052
rect 11701 22043 11759 22049
rect 11790 22040 11796 22052
rect 11848 22080 11854 22092
rect 12452 22080 12480 22120
rect 18325 22083 18383 22089
rect 11848 22052 12480 22080
rect 12728 22052 13032 22080
rect 11848 22040 11854 22052
rect 7285 22015 7343 22021
rect 7285 21981 7297 22015
rect 7331 21981 7343 22015
rect 7285 21975 7343 21981
rect 7377 22015 7435 22021
rect 7377 21981 7389 22015
rect 7423 21981 7435 22015
rect 7377 21975 7435 21981
rect 7561 22015 7619 22021
rect 7561 21981 7573 22015
rect 7607 22012 7619 22015
rect 7742 22012 7748 22024
rect 7607 21984 7748 22012
rect 7607 21981 7619 21984
rect 7561 21975 7619 21981
rect 6730 21904 6736 21956
rect 6788 21944 6794 21956
rect 7392 21944 7420 21975
rect 7742 21972 7748 21984
rect 7800 21972 7806 22024
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 21981 12035 22015
rect 11977 21975 12035 21981
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 12434 22012 12440 22024
rect 12207 21984 12440 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 6788 21916 7420 21944
rect 6788 21904 6794 21916
rect 6362 21836 6368 21888
rect 6420 21836 6426 21888
rect 11992 21876 12020 21975
rect 12434 21972 12440 21984
rect 12492 21972 12498 22024
rect 12526 21972 12532 22024
rect 12584 22012 12590 22024
rect 12728 22021 12756 22052
rect 13004 22024 13032 22052
rect 18325 22049 18337 22083
rect 18371 22080 18383 22083
rect 19426 22080 19432 22092
rect 18371 22052 19432 22080
rect 18371 22049 18383 22052
rect 18325 22043 18383 22049
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 12621 22015 12679 22021
rect 12621 22012 12633 22015
rect 12584 21984 12633 22012
rect 12584 21972 12590 21984
rect 12621 21981 12633 21984
rect 12667 21981 12679 22015
rect 12621 21975 12679 21981
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 21981 12771 22015
rect 12713 21975 12771 21981
rect 12805 22015 12863 22021
rect 12805 21981 12817 22015
rect 12851 21981 12863 22015
rect 12805 21975 12863 21981
rect 12897 22015 12955 22021
rect 12897 21981 12909 22015
rect 12943 21981 12955 22015
rect 12897 21975 12955 21981
rect 12250 21904 12256 21956
rect 12308 21904 12314 21956
rect 12342 21904 12348 21956
rect 12400 21944 12406 21956
rect 12820 21944 12848 21975
rect 12400 21916 12848 21944
rect 12912 21944 12940 21975
rect 12986 21972 12992 22024
rect 13044 21972 13050 22024
rect 17126 21972 17132 22024
rect 17184 22021 17190 22024
rect 17184 21975 17196 22021
rect 17184 21972 17190 21975
rect 17402 21972 17408 22024
rect 17460 22012 17466 22024
rect 18046 22012 18052 22024
rect 17460 21984 18052 22012
rect 17460 21972 17466 21984
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 18509 22015 18567 22021
rect 18509 21981 18521 22015
rect 18555 22012 18567 22015
rect 18598 22012 18604 22024
rect 18555 21984 18604 22012
rect 18555 21981 18567 21984
rect 18509 21975 18567 21981
rect 18598 21972 18604 21984
rect 18656 21972 18662 22024
rect 18782 21972 18788 22024
rect 18840 21972 18846 22024
rect 18966 21972 18972 22024
rect 19024 21972 19030 22024
rect 13814 21944 13820 21956
rect 12912 21916 13820 21944
rect 12400 21904 12406 21916
rect 12912 21876 12940 21916
rect 13814 21904 13820 21916
rect 13872 21944 13878 21956
rect 14642 21944 14648 21956
rect 13872 21916 14648 21944
rect 13872 21904 13878 21916
rect 14642 21904 14648 21916
rect 14700 21904 14706 21956
rect 17954 21904 17960 21956
rect 18012 21944 18018 21956
rect 18877 21947 18935 21953
rect 18877 21944 18889 21947
rect 18012 21916 18889 21944
rect 18012 21904 18018 21916
rect 18877 21913 18889 21916
rect 18923 21913 18935 21947
rect 18877 21907 18935 21913
rect 11992 21848 12940 21876
rect 12986 21836 12992 21888
rect 13044 21876 13050 21888
rect 13173 21879 13231 21885
rect 13173 21876 13185 21879
rect 13044 21848 13185 21876
rect 13044 21836 13050 21848
rect 13173 21845 13185 21848
rect 13219 21845 13231 21879
rect 13173 21839 13231 21845
rect 16025 21879 16083 21885
rect 16025 21845 16037 21879
rect 16071 21876 16083 21879
rect 16574 21876 16580 21888
rect 16071 21848 16580 21876
rect 16071 21845 16083 21848
rect 16025 21839 16083 21845
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 18506 21836 18512 21888
rect 18564 21876 18570 21888
rect 18984 21876 19012 21972
rect 18564 21848 19012 21876
rect 18564 21836 18570 21848
rect 1104 21786 28888 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 28888 21786
rect 1104 21712 28888 21734
rect 12434 21564 12440 21616
rect 12492 21604 12498 21616
rect 12621 21607 12679 21613
rect 12621 21604 12633 21607
rect 12492 21576 12633 21604
rect 12492 21564 12498 21576
rect 12621 21573 12633 21576
rect 12667 21573 12679 21607
rect 12621 21567 12679 21573
rect 12345 21403 12403 21409
rect 12345 21369 12357 21403
rect 12391 21400 12403 21403
rect 12986 21400 12992 21412
rect 12391 21372 12992 21400
rect 12391 21369 12403 21372
rect 12345 21363 12403 21369
rect 12986 21360 12992 21372
rect 13044 21360 13050 21412
rect 12158 21292 12164 21344
rect 12216 21292 12222 21344
rect 1104 21242 28888 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 28888 21242
rect 1104 21168 28888 21190
rect 7006 21088 7012 21140
rect 7064 21128 7070 21140
rect 7190 21128 7196 21140
rect 7064 21100 7196 21128
rect 7064 21088 7070 21100
rect 7190 21088 7196 21100
rect 7248 21128 7254 21140
rect 7561 21131 7619 21137
rect 7561 21128 7573 21131
rect 7248 21100 7573 21128
rect 7248 21088 7254 21100
rect 7561 21097 7573 21100
rect 7607 21097 7619 21131
rect 7561 21091 7619 21097
rect 7006 20884 7012 20936
rect 7064 20884 7070 20936
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 12805 20927 12863 20933
rect 12805 20924 12817 20927
rect 12492 20896 12817 20924
rect 12492 20884 12498 20896
rect 12805 20893 12817 20896
rect 12851 20893 12863 20927
rect 12805 20887 12863 20893
rect 12894 20884 12900 20936
rect 12952 20924 12958 20936
rect 12989 20927 13047 20933
rect 12989 20924 13001 20927
rect 12952 20896 13001 20924
rect 12952 20884 12958 20896
rect 12989 20893 13001 20896
rect 13035 20924 13047 20927
rect 13170 20924 13176 20936
rect 13035 20896 13176 20924
rect 13035 20893 13047 20896
rect 12989 20887 13047 20893
rect 13170 20884 13176 20896
rect 13228 20884 13234 20936
rect 7837 20859 7895 20865
rect 7837 20825 7849 20859
rect 7883 20856 7895 20859
rect 8294 20856 8300 20868
rect 7883 20828 8300 20856
rect 7883 20825 7895 20828
rect 7837 20819 7895 20825
rect 8294 20816 8300 20828
rect 8352 20816 8358 20868
rect 12986 20748 12992 20800
rect 13044 20748 13050 20800
rect 1104 20698 28888 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 28888 20698
rect 1104 20624 28888 20646
rect 16666 20584 16672 20596
rect 9508 20556 16672 20584
rect 9508 20528 9536 20556
rect 16666 20544 16672 20556
rect 16724 20544 16730 20596
rect 9490 20476 9496 20528
rect 9548 20476 9554 20528
rect 13814 20516 13820 20528
rect 12820 20488 13820 20516
rect 5905 20451 5963 20457
rect 5905 20417 5917 20451
rect 5951 20417 5963 20451
rect 5905 20411 5963 20417
rect 6089 20451 6147 20457
rect 6089 20417 6101 20451
rect 6135 20448 6147 20451
rect 6362 20448 6368 20460
rect 6135 20420 6368 20448
rect 6135 20417 6147 20420
rect 6089 20411 6147 20417
rect 5920 20380 5948 20411
rect 6362 20408 6368 20420
rect 6420 20408 6426 20460
rect 12820 20457 12848 20488
rect 13814 20476 13820 20488
rect 13872 20476 13878 20528
rect 14366 20476 14372 20528
rect 14424 20516 14430 20528
rect 17402 20516 17408 20528
rect 14424 20488 17408 20516
rect 14424 20476 14430 20488
rect 14752 20460 14780 20488
rect 17402 20476 17408 20488
rect 17460 20476 17466 20528
rect 12069 20451 12127 20457
rect 12069 20417 12081 20451
rect 12115 20448 12127 20451
rect 12805 20451 12863 20457
rect 12115 20420 12287 20448
rect 12115 20417 12127 20420
rect 12069 20411 12127 20417
rect 7374 20380 7380 20392
rect 5920 20352 7380 20380
rect 7374 20340 7380 20352
rect 7432 20380 7438 20392
rect 8202 20380 8208 20392
rect 7432 20352 8208 20380
rect 7432 20340 7438 20352
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 12158 20340 12164 20392
rect 12216 20340 12222 20392
rect 12259 20380 12287 20420
rect 12805 20417 12817 20451
rect 12851 20417 12863 20451
rect 12805 20411 12863 20417
rect 12894 20408 12900 20460
rect 12952 20408 12958 20460
rect 12986 20408 12992 20460
rect 13044 20408 13050 20460
rect 13078 20408 13084 20460
rect 13136 20448 13142 20460
rect 13173 20451 13231 20457
rect 13173 20448 13185 20451
rect 13136 20420 13185 20448
rect 13136 20408 13142 20420
rect 13173 20417 13185 20420
rect 13219 20448 13231 20451
rect 13262 20448 13268 20460
rect 13219 20420 13268 20448
rect 13219 20417 13231 20420
rect 13173 20411 13231 20417
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 14458 20408 14464 20460
rect 14516 20457 14522 20460
rect 14516 20411 14528 20457
rect 14516 20408 14522 20411
rect 14734 20408 14740 20460
rect 14792 20408 14798 20460
rect 14826 20408 14832 20460
rect 14884 20408 14890 20460
rect 14921 20451 14979 20457
rect 14921 20417 14933 20451
rect 14967 20417 14979 20451
rect 14921 20411 14979 20417
rect 15105 20451 15163 20457
rect 15105 20417 15117 20451
rect 15151 20448 15163 20451
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15151 20420 15853 20448
rect 15151 20417 15163 20420
rect 15105 20411 15163 20417
rect 15841 20417 15853 20420
rect 15887 20448 15899 20451
rect 15930 20448 15936 20460
rect 15887 20420 15936 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 12526 20380 12532 20392
rect 12259 20352 12532 20380
rect 12526 20340 12532 20352
rect 12584 20380 12590 20392
rect 14936 20380 14964 20411
rect 15930 20408 15936 20420
rect 15988 20408 15994 20460
rect 16022 20408 16028 20460
rect 16080 20408 16086 20460
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20448 16175 20451
rect 16298 20448 16304 20460
rect 16163 20420 16304 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 16298 20408 16304 20420
rect 16356 20408 16362 20460
rect 15378 20380 15384 20392
rect 12584 20352 13400 20380
rect 14936 20352 15384 20380
rect 12584 20340 12590 20352
rect 12434 20272 12440 20324
rect 12492 20272 12498 20324
rect 5626 20204 5632 20256
rect 5684 20244 5690 20256
rect 5721 20247 5779 20253
rect 5721 20244 5733 20247
rect 5684 20216 5733 20244
rect 5684 20204 5690 20216
rect 5721 20213 5733 20216
rect 5767 20213 5779 20247
rect 5721 20207 5779 20213
rect 8205 20247 8263 20253
rect 8205 20213 8217 20247
rect 8251 20244 8263 20247
rect 8294 20244 8300 20256
rect 8251 20216 8300 20244
rect 8251 20213 8263 20216
rect 8205 20207 8263 20213
rect 8294 20204 8300 20216
rect 8352 20244 8358 20256
rect 8938 20244 8944 20256
rect 8352 20216 8944 20244
rect 8352 20204 8358 20216
rect 8938 20204 8944 20216
rect 8996 20204 9002 20256
rect 12526 20204 12532 20256
rect 12584 20204 12590 20256
rect 13372 20253 13400 20352
rect 15378 20340 15384 20352
rect 15436 20340 15442 20392
rect 13357 20247 13415 20253
rect 13357 20213 13369 20247
rect 13403 20244 13415 20247
rect 13446 20244 13452 20256
rect 13403 20216 13452 20244
rect 13403 20213 13415 20216
rect 13357 20207 13415 20213
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 14366 20204 14372 20256
rect 14424 20244 14430 20256
rect 15105 20247 15163 20253
rect 15105 20244 15117 20247
rect 14424 20216 15117 20244
rect 14424 20204 14430 20216
rect 15105 20213 15117 20216
rect 15151 20213 15163 20247
rect 15105 20207 15163 20213
rect 15838 20204 15844 20256
rect 15896 20204 15902 20256
rect 1104 20154 28888 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 28888 20154
rect 1104 20080 28888 20102
rect 6822 20000 6828 20052
rect 6880 20000 6886 20052
rect 13170 20000 13176 20052
rect 13228 20040 13234 20052
rect 14185 20043 14243 20049
rect 14185 20040 14197 20043
rect 13228 20012 14197 20040
rect 13228 20000 13234 20012
rect 14185 20009 14197 20012
rect 14231 20009 14243 20043
rect 14185 20003 14243 20009
rect 13814 19932 13820 19984
rect 13872 19932 13878 19984
rect 14200 19972 14228 20003
rect 14458 20000 14464 20052
rect 14516 20040 14522 20052
rect 14553 20043 14611 20049
rect 14553 20040 14565 20043
rect 14516 20012 14565 20040
rect 14516 20000 14522 20012
rect 14553 20009 14565 20012
rect 14599 20009 14611 20043
rect 14553 20003 14611 20009
rect 16298 20000 16304 20052
rect 16356 20040 16362 20052
rect 16669 20043 16727 20049
rect 16669 20040 16681 20043
rect 16356 20012 16681 20040
rect 16356 20000 16362 20012
rect 16669 20009 16681 20012
rect 16715 20009 16727 20043
rect 16669 20003 16727 20009
rect 14826 19972 14832 19984
rect 14200 19944 14832 19972
rect 14826 19932 14832 19944
rect 14884 19932 14890 19984
rect 5350 19864 5356 19916
rect 5408 19904 5414 19916
rect 5445 19907 5503 19913
rect 5445 19904 5457 19907
rect 5408 19876 5457 19904
rect 5408 19864 5414 19876
rect 5445 19873 5457 19876
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 13446 19864 13452 19916
rect 13504 19904 13510 19916
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 13504 19876 14105 19904
rect 13504 19864 13510 19876
rect 14093 19873 14105 19876
rect 14139 19904 14151 19907
rect 14139 19876 14504 19904
rect 14139 19873 14151 19876
rect 14093 19867 14151 19873
rect 6178 19796 6184 19848
rect 6236 19836 6242 19848
rect 6730 19836 6736 19848
rect 6236 19808 6736 19836
rect 6236 19796 6242 19808
rect 6730 19796 6736 19808
rect 6788 19836 6794 19848
rect 7469 19839 7527 19845
rect 7469 19836 7481 19839
rect 6788 19808 7481 19836
rect 6788 19796 6794 19808
rect 7469 19805 7481 19808
rect 7515 19805 7527 19839
rect 7469 19799 7527 19805
rect 8938 19796 8944 19848
rect 8996 19836 9002 19848
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 8996 19808 12449 19836
rect 8996 19796 9002 19808
rect 12437 19805 12449 19808
rect 12483 19805 12495 19839
rect 12437 19799 12495 19805
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 12693 19839 12751 19845
rect 12693 19836 12705 19839
rect 12584 19808 12705 19836
rect 12584 19796 12590 19808
rect 12693 19805 12705 19808
rect 12739 19805 12751 19839
rect 12693 19799 12751 19805
rect 14366 19796 14372 19848
rect 14424 19796 14430 19848
rect 14476 19836 14504 19876
rect 14734 19864 14740 19916
rect 14792 19904 14798 19916
rect 15289 19907 15347 19913
rect 15289 19904 15301 19907
rect 14792 19876 15301 19904
rect 14792 19864 14798 19876
rect 15289 19873 15301 19876
rect 15335 19873 15347 19907
rect 16684 19904 16712 20003
rect 17313 19907 17371 19913
rect 17313 19904 17325 19907
rect 16684 19876 17325 19904
rect 15289 19867 15347 19873
rect 17313 19873 17325 19876
rect 17359 19873 17371 19907
rect 17313 19867 17371 19873
rect 15378 19836 15384 19848
rect 14476 19808 15384 19836
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 28534 19796 28540 19848
rect 28592 19796 28598 19848
rect 5712 19771 5770 19777
rect 5712 19737 5724 19771
rect 5758 19768 5770 19771
rect 6362 19768 6368 19780
rect 5758 19740 6368 19768
rect 5758 19737 5770 19740
rect 5712 19731 5770 19737
rect 6362 19728 6368 19740
rect 6420 19728 6426 19780
rect 15556 19771 15614 19777
rect 15556 19737 15568 19771
rect 15602 19768 15614 19771
rect 15654 19768 15660 19780
rect 15602 19740 15660 19768
rect 15602 19737 15614 19740
rect 15556 19731 15614 19737
rect 15654 19728 15660 19740
rect 15712 19728 15718 19780
rect 6914 19660 6920 19712
rect 6972 19660 6978 19712
rect 16758 19660 16764 19712
rect 16816 19660 16822 19712
rect 1104 19610 28888 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 28888 19610
rect 1104 19536 28888 19558
rect 6178 19456 6184 19508
rect 6236 19456 6242 19508
rect 6362 19456 6368 19508
rect 6420 19456 6426 19508
rect 7374 19456 7380 19508
rect 7432 19456 7438 19508
rect 15654 19456 15660 19508
rect 15712 19456 15718 19508
rect 5350 19428 5356 19440
rect 4816 19400 5356 19428
rect 4816 19369 4844 19400
rect 5350 19388 5356 19400
rect 5408 19388 5414 19440
rect 6825 19431 6883 19437
rect 6825 19428 6837 19431
rect 5920 19400 6837 19428
rect 4801 19363 4859 19369
rect 4801 19329 4813 19363
rect 4847 19329 4859 19363
rect 4801 19323 4859 19329
rect 5068 19363 5126 19369
rect 5068 19329 5080 19363
rect 5114 19360 5126 19363
rect 5920 19360 5948 19400
rect 6825 19397 6837 19400
rect 6871 19397 6883 19431
rect 6825 19391 6883 19397
rect 5114 19332 5948 19360
rect 6549 19363 6607 19369
rect 5114 19329 5126 19332
rect 5068 19323 5126 19329
rect 6549 19329 6561 19363
rect 6595 19360 6607 19363
rect 7009 19363 7067 19369
rect 7009 19360 7021 19363
rect 6595 19332 7021 19360
rect 6595 19329 6607 19332
rect 6549 19323 6607 19329
rect 7009 19329 7021 19332
rect 7055 19360 7067 19363
rect 7392 19360 7420 19456
rect 16758 19428 16764 19440
rect 16040 19400 16764 19428
rect 7055 19332 7420 19360
rect 7469 19363 7527 19369
rect 7055 19329 7067 19332
rect 7009 19323 7067 19329
rect 7469 19329 7481 19363
rect 7515 19360 7527 19363
rect 8846 19360 8852 19372
rect 7515 19332 8852 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 15838 19320 15844 19372
rect 15896 19320 15902 19372
rect 16040 19369 16068 19400
rect 16758 19388 16764 19400
rect 16816 19388 16822 19440
rect 16025 19363 16083 19369
rect 16025 19329 16037 19363
rect 16071 19329 16083 19363
rect 16025 19323 16083 19329
rect 16114 19320 16120 19372
rect 16172 19320 16178 19372
rect 16666 19320 16672 19372
rect 16724 19360 16730 19372
rect 17954 19360 17960 19372
rect 16724 19332 17960 19360
rect 16724 19320 16730 19332
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 6733 19295 6791 19301
rect 6733 19261 6745 19295
rect 6779 19292 6791 19295
rect 6914 19292 6920 19304
rect 6779 19264 6920 19292
rect 6779 19261 6791 19264
rect 6733 19255 6791 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 7190 19252 7196 19304
rect 7248 19252 7254 19304
rect 9585 19295 9643 19301
rect 9585 19261 9597 19295
rect 9631 19292 9643 19295
rect 9766 19292 9772 19304
rect 9631 19264 9772 19292
rect 9631 19261 9643 19264
rect 9585 19255 9643 19261
rect 9766 19252 9772 19264
rect 9824 19252 9830 19304
rect 8754 19116 8760 19168
rect 8812 19156 8818 19168
rect 8941 19159 8999 19165
rect 8941 19156 8953 19159
rect 8812 19128 8953 19156
rect 8812 19116 8818 19128
rect 8941 19125 8953 19128
rect 8987 19125 8999 19159
rect 8941 19119 8999 19125
rect 1104 19066 28888 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 28888 19066
rect 1104 18992 28888 19014
rect 6733 18955 6791 18961
rect 6733 18921 6745 18955
rect 6779 18952 6791 18955
rect 7006 18952 7012 18964
rect 6779 18924 7012 18952
rect 6779 18921 6791 18924
rect 6733 18915 6791 18921
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 22094 18844 22100 18896
rect 22152 18884 22158 18896
rect 23385 18887 23443 18893
rect 23385 18884 23397 18887
rect 22152 18856 23397 18884
rect 22152 18844 22158 18856
rect 23385 18853 23397 18856
rect 23431 18853 23443 18887
rect 23385 18847 23443 18853
rect 5350 18776 5356 18828
rect 5408 18776 5414 18828
rect 8938 18776 8944 18828
rect 8996 18776 9002 18828
rect 21082 18776 21088 18828
rect 21140 18816 21146 18828
rect 21361 18819 21419 18825
rect 21361 18816 21373 18819
rect 21140 18788 21373 18816
rect 21140 18776 21146 18788
rect 21361 18785 21373 18788
rect 21407 18785 21419 18819
rect 21361 18779 21419 18785
rect 21468 18788 23060 18816
rect 21468 18760 21496 18788
rect 5626 18757 5632 18760
rect 5620 18748 5632 18757
rect 5587 18720 5632 18748
rect 5620 18711 5632 18720
rect 5626 18708 5632 18711
rect 5684 18708 5690 18760
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 19300 18720 19533 18748
rect 19300 18708 19306 18720
rect 19521 18717 19533 18720
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 20993 18751 21051 18757
rect 20993 18748 21005 18751
rect 20956 18720 21005 18748
rect 20956 18708 20962 18720
rect 20993 18717 21005 18720
rect 21039 18717 21051 18751
rect 20993 18711 21051 18717
rect 21174 18708 21180 18760
rect 21232 18708 21238 18760
rect 21450 18708 21456 18760
rect 21508 18708 21514 18760
rect 21637 18751 21695 18757
rect 21637 18717 21649 18751
rect 21683 18748 21695 18751
rect 22094 18748 22100 18760
rect 21683 18720 22100 18748
rect 21683 18717 21695 18720
rect 21637 18711 21695 18717
rect 22094 18708 22100 18720
rect 22152 18708 22158 18760
rect 23032 18757 23060 18788
rect 22925 18751 22983 18757
rect 22925 18717 22937 18751
rect 22971 18717 22983 18751
rect 22925 18711 22983 18717
rect 23017 18751 23075 18757
rect 23017 18717 23029 18751
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 23569 18751 23627 18757
rect 23569 18717 23581 18751
rect 23615 18748 23627 18751
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 23615 18720 23765 18748
rect 23615 18717 23627 18720
rect 23569 18711 23627 18717
rect 23753 18717 23765 18720
rect 23799 18717 23811 18751
rect 23753 18711 23811 18717
rect 9030 18640 9036 18692
rect 9088 18680 9094 18692
rect 9186 18683 9244 18689
rect 9186 18680 9198 18683
rect 9088 18652 9198 18680
rect 9088 18640 9094 18652
rect 9186 18649 9198 18652
rect 9232 18649 9244 18683
rect 9186 18643 9244 18649
rect 19610 18640 19616 18692
rect 19668 18680 19674 18692
rect 19766 18683 19824 18689
rect 19766 18680 19778 18683
rect 19668 18652 19778 18680
rect 19668 18640 19674 18652
rect 19766 18649 19778 18652
rect 19812 18649 19824 18683
rect 19766 18643 19824 18649
rect 20714 18640 20720 18692
rect 20772 18680 20778 18692
rect 21545 18683 21603 18689
rect 21545 18680 21557 18683
rect 20772 18652 21557 18680
rect 20772 18640 20778 18652
rect 21545 18649 21557 18652
rect 21591 18649 21603 18683
rect 22940 18680 22968 18711
rect 23658 18680 23664 18692
rect 22940 18652 23664 18680
rect 21545 18643 21603 18649
rect 23658 18640 23664 18652
rect 23716 18640 23722 18692
rect 23768 18680 23796 18711
rect 23934 18708 23940 18760
rect 23992 18708 23998 18760
rect 25498 18680 25504 18692
rect 23768 18652 25504 18680
rect 25498 18640 25504 18652
rect 25556 18680 25562 18692
rect 27522 18680 27528 18692
rect 25556 18652 27528 18680
rect 25556 18640 25562 18652
rect 27522 18640 27528 18652
rect 27580 18640 27586 18692
rect 10318 18572 10324 18624
rect 10376 18572 10382 18624
rect 20901 18615 20959 18621
rect 20901 18581 20913 18615
rect 20947 18612 20959 18615
rect 21082 18612 21088 18624
rect 20947 18584 21088 18612
rect 20947 18581 20959 18584
rect 20901 18575 20959 18581
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 23106 18572 23112 18624
rect 23164 18612 23170 18624
rect 23201 18615 23259 18621
rect 23201 18612 23213 18615
rect 23164 18584 23213 18612
rect 23164 18572 23170 18584
rect 23201 18581 23213 18584
rect 23247 18581 23259 18615
rect 23201 18575 23259 18581
rect 23474 18572 23480 18624
rect 23532 18612 23538 18624
rect 23845 18615 23903 18621
rect 23845 18612 23857 18615
rect 23532 18584 23857 18612
rect 23532 18572 23538 18584
rect 23845 18581 23857 18584
rect 23891 18581 23903 18615
rect 23845 18575 23903 18581
rect 1104 18522 28888 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 28888 18522
rect 1104 18448 28888 18470
rect 9030 18368 9036 18420
rect 9088 18368 9094 18420
rect 23385 18411 23443 18417
rect 23385 18377 23397 18411
rect 23431 18408 23443 18411
rect 23658 18408 23664 18420
rect 23431 18380 23664 18408
rect 23431 18377 23443 18380
rect 23385 18371 23443 18377
rect 23658 18368 23664 18380
rect 23716 18368 23722 18420
rect 13170 18340 13176 18352
rect 9784 18312 13176 18340
rect 8754 18232 8760 18284
rect 8812 18232 8818 18284
rect 8846 18232 8852 18284
rect 8904 18281 8910 18284
rect 8904 18275 8927 18281
rect 8915 18272 8927 18275
rect 9784 18272 9812 18312
rect 13170 18300 13176 18312
rect 13228 18300 13234 18352
rect 20180 18312 24992 18340
rect 8915 18244 9812 18272
rect 8915 18241 8927 18244
rect 8904 18235 8927 18241
rect 8904 18232 8910 18235
rect 9858 18232 9864 18284
rect 9916 18272 9922 18284
rect 10238 18275 10296 18281
rect 10238 18272 10250 18275
rect 9916 18244 10250 18272
rect 9916 18232 9922 18244
rect 10238 18241 10250 18244
rect 10284 18241 10296 18275
rect 10238 18235 10296 18241
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18241 15255 18275
rect 15197 18235 15255 18241
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18272 15439 18275
rect 15749 18275 15807 18281
rect 15749 18272 15761 18275
rect 15427 18244 15761 18272
rect 15427 18241 15439 18244
rect 15381 18235 15439 18241
rect 15749 18241 15761 18244
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 10505 18207 10563 18213
rect 10505 18173 10517 18207
rect 10551 18204 10563 18207
rect 11330 18204 11336 18216
rect 10551 18176 11336 18204
rect 10551 18173 10563 18176
rect 10505 18167 10563 18173
rect 11330 18164 11336 18176
rect 11388 18164 11394 18216
rect 15212 18204 15240 18235
rect 16114 18232 16120 18284
rect 16172 18272 16178 18284
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 16172 18244 16313 18272
rect 16172 18232 16178 18244
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 16301 18235 16359 18241
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18690 18272 18696 18284
rect 18012 18244 18696 18272
rect 18012 18232 18018 18244
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 20180 18281 20208 18312
rect 20438 18281 20444 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 19300 18244 20177 18272
rect 19300 18232 19306 18244
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 20432 18235 20444 18281
rect 20438 18232 20444 18235
rect 20496 18232 20502 18284
rect 22020 18281 22048 18312
rect 22278 18281 22284 18284
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22272 18235 22284 18281
rect 22278 18232 22284 18235
rect 22336 18232 22342 18284
rect 23492 18281 23520 18312
rect 23750 18281 23756 18284
rect 23477 18275 23535 18281
rect 23477 18241 23489 18275
rect 23523 18241 23535 18275
rect 23477 18235 23535 18241
rect 23744 18235 23756 18281
rect 23750 18232 23756 18235
rect 23808 18232 23814 18284
rect 15930 18204 15936 18216
rect 15212 18176 15936 18204
rect 15930 18164 15936 18176
rect 15988 18204 15994 18216
rect 18506 18204 18512 18216
rect 15988 18176 18512 18204
rect 15988 18164 15994 18176
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 24964 18213 24992 18312
rect 25222 18281 25228 18284
rect 25216 18235 25228 18281
rect 25222 18232 25228 18235
rect 25280 18232 25286 18284
rect 24949 18207 25007 18213
rect 24949 18173 24961 18207
rect 24995 18173 25007 18207
rect 24949 18167 25007 18173
rect 9125 18071 9183 18077
rect 9125 18037 9137 18071
rect 9171 18068 9183 18071
rect 9766 18068 9772 18080
rect 9171 18040 9772 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9766 18028 9772 18040
rect 9824 18068 9830 18080
rect 10502 18068 10508 18080
rect 9824 18040 10508 18068
rect 9824 18028 9830 18040
rect 10502 18028 10508 18040
rect 10560 18028 10566 18080
rect 15194 18028 15200 18080
rect 15252 18028 15258 18080
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 19242 18068 19248 18080
rect 18380 18040 19248 18068
rect 18380 18028 18386 18040
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 21542 18028 21548 18080
rect 21600 18028 21606 18080
rect 24854 18028 24860 18080
rect 24912 18028 24918 18080
rect 24964 18068 24992 18167
rect 26234 18068 26240 18080
rect 24964 18040 26240 18068
rect 26234 18028 26240 18040
rect 26292 18028 26298 18080
rect 26329 18071 26387 18077
rect 26329 18037 26341 18071
rect 26375 18068 26387 18071
rect 26510 18068 26516 18080
rect 26375 18040 26516 18068
rect 26375 18037 26387 18040
rect 26329 18031 26387 18037
rect 26510 18028 26516 18040
rect 26568 18028 26574 18080
rect 1104 17978 28888 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 28888 17978
rect 1104 17904 28888 17926
rect 16025 17867 16083 17873
rect 16025 17833 16037 17867
rect 16071 17864 16083 17867
rect 16114 17864 16120 17876
rect 16071 17836 16120 17864
rect 16071 17833 16083 17836
rect 16025 17827 16083 17833
rect 16114 17824 16120 17836
rect 16172 17824 16178 17876
rect 19610 17824 19616 17876
rect 19668 17824 19674 17876
rect 22278 17824 22284 17876
rect 22336 17864 22342 17876
rect 22373 17867 22431 17873
rect 22373 17864 22385 17867
rect 22336 17836 22385 17864
rect 22336 17824 22342 17836
rect 22373 17833 22385 17836
rect 22419 17833 22431 17867
rect 22373 17827 22431 17833
rect 23845 17867 23903 17873
rect 23845 17833 23857 17867
rect 23891 17864 23903 17867
rect 23934 17864 23940 17876
rect 23891 17836 23940 17864
rect 23891 17833 23903 17836
rect 23845 17827 23903 17833
rect 23934 17824 23940 17836
rect 23992 17824 23998 17876
rect 24026 17824 24032 17876
rect 24084 17824 24090 17876
rect 25133 17867 25191 17873
rect 25133 17833 25145 17867
rect 25179 17864 25191 17867
rect 25222 17864 25228 17876
rect 25179 17836 25228 17864
rect 25179 17833 25191 17836
rect 25133 17827 25191 17833
rect 25222 17824 25228 17836
rect 25280 17824 25286 17876
rect 19981 17799 20039 17805
rect 19981 17796 19993 17799
rect 18800 17768 19993 17796
rect 10137 17663 10195 17669
rect 10137 17629 10149 17663
rect 10183 17660 10195 17663
rect 10226 17660 10232 17672
rect 10183 17632 10232 17660
rect 10183 17629 10195 17632
rect 10137 17623 10195 17629
rect 10226 17620 10232 17632
rect 10284 17620 10290 17672
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 10778 17660 10784 17672
rect 10367 17632 10784 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17660 14703 17663
rect 14734 17660 14740 17672
rect 14691 17632 14740 17660
rect 14691 17629 14703 17632
rect 14645 17623 14703 17629
rect 14734 17620 14740 17632
rect 14792 17660 14798 17672
rect 18322 17660 18328 17672
rect 14792 17632 18328 17660
rect 14792 17620 14798 17632
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 18414 17620 18420 17672
rect 18472 17660 18478 17672
rect 18800 17669 18828 17768
rect 19981 17765 19993 17768
rect 20027 17796 20039 17799
rect 21174 17796 21180 17808
rect 20027 17768 21180 17796
rect 20027 17765 20039 17768
rect 19981 17759 20039 17765
rect 21174 17756 21180 17768
rect 21232 17756 21238 17808
rect 21450 17756 21456 17808
rect 21508 17796 21514 17808
rect 22741 17799 22799 17805
rect 22741 17796 22753 17799
rect 21508 17768 22753 17796
rect 21508 17756 21514 17768
rect 22741 17765 22753 17768
rect 22787 17765 22799 17799
rect 23952 17796 23980 17824
rect 24762 17796 24768 17808
rect 23952 17768 24768 17796
rect 22741 17759 22799 17765
rect 20257 17731 20315 17737
rect 20257 17728 20269 17731
rect 19812 17700 20269 17728
rect 18693 17663 18751 17669
rect 18693 17660 18705 17663
rect 18472 17632 18705 17660
rect 18472 17620 18478 17632
rect 18693 17629 18705 17632
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 18785 17663 18843 17669
rect 18785 17629 18797 17663
rect 18831 17660 18843 17663
rect 18874 17660 18880 17672
rect 18831 17632 18880 17660
rect 18831 17629 18843 17632
rect 18785 17623 18843 17629
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 19812 17669 19840 17700
rect 20257 17697 20269 17700
rect 20303 17697 20315 17731
rect 20257 17691 20315 17697
rect 20806 17688 20812 17740
rect 20864 17728 20870 17740
rect 21542 17728 21548 17740
rect 20864 17700 21548 17728
rect 20864 17688 20870 17700
rect 21542 17688 21548 17700
rect 21600 17728 21606 17740
rect 21821 17731 21879 17737
rect 21821 17728 21833 17731
rect 21600 17700 21833 17728
rect 21600 17688 21606 17700
rect 21821 17697 21833 17700
rect 21867 17697 21879 17731
rect 21821 17691 21879 17697
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17629 20131 17663
rect 20073 17623 20131 17629
rect 14912 17595 14970 17601
rect 14912 17561 14924 17595
rect 14958 17592 14970 17595
rect 15194 17592 15200 17604
rect 14958 17564 15200 17592
rect 14958 17561 14970 17564
rect 14912 17555 14970 17561
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 18506 17552 18512 17604
rect 18564 17592 18570 17604
rect 20088 17592 20116 17623
rect 20162 17620 20168 17672
rect 20220 17620 20226 17672
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17660 20407 17663
rect 20898 17660 20904 17672
rect 20395 17632 20904 17660
rect 20395 17629 20407 17632
rect 20349 17623 20407 17629
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 21082 17620 21088 17672
rect 21140 17620 21146 17672
rect 22554 17620 22560 17672
rect 22612 17620 22618 17672
rect 20533 17595 20591 17601
rect 20533 17592 20545 17595
rect 18564 17564 18920 17592
rect 20088 17564 20545 17592
rect 18564 17552 18570 17564
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 9953 17527 10011 17533
rect 9953 17524 9965 17527
rect 9916 17496 9965 17524
rect 9916 17484 9922 17496
rect 9953 17493 9965 17496
rect 9999 17493 10011 17527
rect 9953 17487 10011 17493
rect 18782 17484 18788 17536
rect 18840 17484 18846 17536
rect 18892 17524 18920 17564
rect 20533 17561 20545 17564
rect 20579 17561 20591 17595
rect 22094 17592 22100 17604
rect 20533 17555 20591 17561
rect 20640 17564 22100 17592
rect 20162 17524 20168 17536
rect 18892 17496 20168 17524
rect 20162 17484 20168 17496
rect 20220 17524 20226 17536
rect 20640 17524 20668 17564
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 22756 17592 22784 17759
rect 24762 17756 24768 17768
rect 24820 17796 24826 17808
rect 25501 17799 25559 17805
rect 25501 17796 25513 17799
rect 24820 17768 25513 17796
rect 24820 17756 24826 17768
rect 25501 17765 25513 17768
rect 25547 17765 25559 17799
rect 25501 17759 25559 17765
rect 23658 17688 23664 17740
rect 23716 17728 23722 17740
rect 24026 17728 24032 17740
rect 23716 17700 24032 17728
rect 23716 17688 23722 17700
rect 24026 17688 24032 17700
rect 24084 17688 24090 17740
rect 25593 17731 25651 17737
rect 25593 17697 25605 17731
rect 25639 17728 25651 17731
rect 25866 17728 25872 17740
rect 25639 17700 25872 17728
rect 25639 17697 25651 17700
rect 25593 17691 25651 17697
rect 25866 17688 25872 17700
rect 25924 17728 25930 17740
rect 26697 17731 26755 17737
rect 26697 17728 26709 17731
rect 25924 17700 26709 17728
rect 25924 17688 25930 17700
rect 26697 17697 26709 17700
rect 26743 17697 26755 17731
rect 26697 17691 26755 17697
rect 22833 17663 22891 17669
rect 22833 17629 22845 17663
rect 22879 17660 22891 17663
rect 23109 17663 23167 17669
rect 23109 17660 23121 17663
rect 22879 17632 23121 17660
rect 22879 17629 22891 17632
rect 22833 17623 22891 17629
rect 23109 17629 23121 17632
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 24949 17663 25007 17669
rect 24949 17629 24961 17663
rect 24995 17629 25007 17663
rect 24949 17623 25007 17629
rect 25317 17663 25375 17669
rect 25317 17629 25329 17663
rect 25363 17660 25375 17663
rect 25406 17660 25412 17672
rect 25363 17632 25412 17660
rect 25363 17629 25375 17632
rect 25317 17623 25375 17629
rect 23997 17595 24055 17601
rect 23997 17592 24009 17595
rect 22756 17564 24009 17592
rect 23997 17561 24009 17564
rect 24043 17561 24055 17595
rect 23997 17555 24055 17561
rect 24213 17595 24271 17601
rect 24213 17561 24225 17595
rect 24259 17592 24271 17595
rect 24302 17592 24308 17604
rect 24259 17564 24308 17592
rect 24259 17561 24271 17564
rect 24213 17555 24271 17561
rect 24302 17552 24308 17564
rect 24360 17592 24366 17604
rect 24854 17592 24860 17604
rect 24360 17564 24860 17592
rect 24360 17552 24366 17564
rect 24854 17552 24860 17564
rect 24912 17592 24918 17604
rect 24964 17592 24992 17623
rect 25406 17620 25412 17632
rect 25464 17620 25470 17672
rect 26510 17620 26516 17672
rect 26568 17660 26574 17672
rect 27249 17663 27307 17669
rect 27249 17660 27261 17663
rect 26568 17632 27261 17660
rect 26568 17620 26574 17632
rect 27249 17629 27261 17632
rect 27295 17629 27307 17663
rect 27249 17623 27307 17629
rect 24912 17564 24992 17592
rect 24912 17552 24918 17564
rect 20220 17496 20668 17524
rect 20220 17484 20226 17496
rect 20990 17484 20996 17536
rect 21048 17524 21054 17536
rect 21269 17527 21327 17533
rect 21269 17524 21281 17527
rect 21048 17496 21281 17524
rect 21048 17484 21054 17496
rect 21269 17493 21281 17496
rect 21315 17493 21327 17527
rect 21269 17487 21327 17493
rect 24394 17484 24400 17536
rect 24452 17484 24458 17536
rect 25590 17484 25596 17536
rect 25648 17524 25654 17536
rect 25961 17527 26019 17533
rect 25961 17524 25973 17527
rect 25648 17496 25973 17524
rect 25648 17484 25654 17496
rect 25961 17493 25973 17496
rect 26007 17493 26019 17527
rect 25961 17487 26019 17493
rect 1104 17434 28888 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 28888 17434
rect 1104 17360 28888 17382
rect 20438 17280 20444 17332
rect 20496 17320 20502 17332
rect 20533 17323 20591 17329
rect 20533 17320 20545 17323
rect 20496 17292 20545 17320
rect 20496 17280 20502 17292
rect 20533 17289 20545 17292
rect 20579 17289 20591 17323
rect 20533 17283 20591 17289
rect 21174 17280 21180 17332
rect 21232 17320 21238 17332
rect 21285 17323 21343 17329
rect 21285 17320 21297 17323
rect 21232 17292 21297 17320
rect 21232 17280 21238 17292
rect 21285 17289 21297 17292
rect 21331 17289 21343 17323
rect 21285 17283 21343 17289
rect 21450 17280 21456 17332
rect 21508 17280 21514 17332
rect 22554 17280 22560 17332
rect 22612 17320 22618 17332
rect 23017 17323 23075 17329
rect 23017 17320 23029 17323
rect 22612 17292 23029 17320
rect 22612 17280 22618 17292
rect 23017 17289 23029 17292
rect 23063 17289 23075 17323
rect 23017 17283 23075 17289
rect 23661 17323 23719 17329
rect 23661 17289 23673 17323
rect 23707 17320 23719 17323
rect 23750 17320 23756 17332
rect 23707 17292 23756 17320
rect 23707 17289 23719 17292
rect 23661 17283 23719 17289
rect 23750 17280 23756 17292
rect 23808 17280 23814 17332
rect 25590 17280 25596 17332
rect 25648 17280 25654 17332
rect 10226 17212 10232 17264
rect 10284 17252 10290 17264
rect 11514 17252 11520 17264
rect 10284 17224 11520 17252
rect 10284 17212 10290 17224
rect 11514 17212 11520 17224
rect 11572 17212 11578 17264
rect 18592 17255 18650 17261
rect 18592 17221 18604 17255
rect 18638 17252 18650 17255
rect 18782 17252 18788 17264
rect 18638 17224 18788 17252
rect 18638 17221 18650 17224
rect 18592 17215 18650 17221
rect 18782 17212 18788 17224
rect 18840 17212 18846 17264
rect 20806 17212 20812 17264
rect 20864 17252 20870 17264
rect 21085 17255 21143 17261
rect 21085 17252 21097 17255
rect 20864 17224 21097 17252
rect 20864 17212 20870 17224
rect 21085 17221 21097 17224
rect 21131 17221 21143 17255
rect 24394 17252 24400 17264
rect 21085 17215 21143 17221
rect 23216 17224 24400 17252
rect 11077 17187 11135 17193
rect 11077 17153 11089 17187
rect 11123 17184 11135 17187
rect 11238 17184 11244 17196
rect 11123 17156 11244 17184
rect 11123 17153 11135 17156
rect 11077 17147 11135 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 11330 17144 11336 17196
rect 11388 17144 11394 17196
rect 16945 17187 17003 17193
rect 16945 17153 16957 17187
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17184 17187 17187
rect 17589 17187 17647 17193
rect 17589 17184 17601 17187
rect 17175 17156 17601 17184
rect 17175 17153 17187 17156
rect 17129 17147 17187 17153
rect 17589 17153 17601 17156
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 16960 17116 16988 17147
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 20714 17144 20720 17196
rect 20772 17144 20778 17196
rect 20898 17144 20904 17196
rect 20956 17144 20962 17196
rect 20990 17144 20996 17196
rect 21048 17144 21054 17196
rect 22094 17144 22100 17196
rect 22152 17184 22158 17196
rect 22925 17187 22983 17193
rect 22925 17184 22937 17187
rect 22152 17156 22937 17184
rect 22152 17144 22158 17156
rect 22925 17153 22937 17156
rect 22971 17153 22983 17187
rect 22925 17147 22983 17153
rect 23106 17144 23112 17196
rect 23164 17144 23170 17196
rect 23216 17193 23244 17224
rect 24394 17212 24400 17224
rect 24452 17212 24458 17264
rect 24762 17212 24768 17264
rect 24820 17252 24826 17264
rect 24820 17224 25728 17252
rect 24820 17212 24826 17224
rect 23201 17187 23259 17193
rect 23201 17153 23213 17187
rect 23247 17153 23259 17187
rect 23201 17147 23259 17153
rect 23474 17144 23480 17196
rect 23532 17144 23538 17196
rect 25409 17187 25467 17193
rect 25409 17153 25421 17187
rect 25455 17184 25467 17187
rect 25498 17184 25504 17196
rect 25455 17156 25504 17184
rect 25455 17153 25467 17156
rect 25409 17147 25467 17153
rect 25498 17144 25504 17156
rect 25556 17144 25562 17196
rect 25700 17193 25728 17224
rect 25685 17187 25743 17193
rect 25685 17153 25697 17187
rect 25731 17153 25743 17187
rect 25685 17147 25743 17153
rect 18138 17116 18144 17128
rect 16960 17088 18144 17116
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 18230 17076 18236 17128
rect 18288 17076 18294 17128
rect 20349 17119 20407 17125
rect 20349 17116 20361 17119
rect 19720 17088 20361 17116
rect 19720 17060 19748 17088
rect 20349 17085 20361 17088
rect 20395 17085 20407 17119
rect 23124 17116 23152 17144
rect 23293 17119 23351 17125
rect 23293 17116 23305 17119
rect 23124 17088 23305 17116
rect 20349 17079 20407 17085
rect 23293 17085 23305 17088
rect 23339 17085 23351 17119
rect 23293 17079 23351 17085
rect 19702 17008 19708 17060
rect 19760 17008 19766 17060
rect 25406 17008 25412 17060
rect 25464 17008 25470 17060
rect 9950 16940 9956 16992
rect 10008 16940 10014 16992
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 12158 16980 12164 16992
rect 11204 16952 12164 16980
rect 11204 16940 11210 16952
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 16850 16940 16856 16992
rect 16908 16980 16914 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16908 16952 16957 16980
rect 16908 16940 16914 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 19794 16940 19800 16992
rect 19852 16940 19858 16992
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 21082 16980 21088 16992
rect 20680 16952 21088 16980
rect 20680 16940 20686 16952
rect 21082 16940 21088 16952
rect 21140 16980 21146 16992
rect 21269 16983 21327 16989
rect 21269 16980 21281 16983
rect 21140 16952 21281 16980
rect 21140 16940 21146 16952
rect 21269 16949 21281 16952
rect 21315 16949 21327 16983
rect 21269 16943 21327 16949
rect 1104 16890 28888 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 28888 16890
rect 1104 16816 28888 16838
rect 9309 16779 9367 16785
rect 9309 16745 9321 16779
rect 9355 16776 9367 16779
rect 9355 16748 11192 16776
rect 9355 16745 9367 16748
rect 9309 16739 9367 16745
rect 9950 16668 9956 16720
rect 10008 16708 10014 16720
rect 10008 16680 10180 16708
rect 10008 16668 10014 16680
rect 10152 16649 10180 16680
rect 10778 16668 10784 16720
rect 10836 16668 10842 16720
rect 11164 16708 11192 16748
rect 11238 16736 11244 16788
rect 11296 16776 11302 16788
rect 11517 16779 11575 16785
rect 11517 16776 11529 16779
rect 11296 16748 11529 16776
rect 11296 16736 11302 16748
rect 11517 16745 11529 16748
rect 11563 16745 11575 16779
rect 11517 16739 11575 16745
rect 12158 16736 12164 16788
rect 12216 16736 12222 16788
rect 18322 16776 18328 16788
rect 16592 16748 18328 16776
rect 11164 16680 11376 16708
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16640 9551 16643
rect 10137 16643 10195 16649
rect 9539 16612 10088 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 5534 16532 5540 16584
rect 5592 16572 5598 16584
rect 6273 16575 6331 16581
rect 6273 16572 6285 16575
rect 5592 16544 6285 16572
rect 5592 16532 5598 16544
rect 6273 16541 6285 16544
rect 6319 16572 6331 16575
rect 7650 16572 7656 16584
rect 6319 16544 7656 16572
rect 6319 16541 6331 16544
rect 6273 16535 6331 16541
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 7745 16575 7803 16581
rect 7745 16541 7757 16575
rect 7791 16572 7803 16575
rect 8294 16572 8300 16584
rect 7791 16544 8300 16572
rect 7791 16541 7803 16544
rect 7745 16535 7803 16541
rect 8294 16532 8300 16544
rect 8352 16572 8358 16584
rect 9585 16575 9643 16581
rect 9585 16572 9597 16575
rect 8352 16544 9597 16572
rect 8352 16532 8358 16544
rect 9585 16541 9597 16544
rect 9631 16541 9643 16575
rect 9585 16535 9643 16541
rect 9858 16532 9864 16584
rect 9916 16532 9922 16584
rect 9950 16532 9956 16584
rect 10008 16532 10014 16584
rect 10060 16572 10088 16612
rect 10137 16609 10149 16643
rect 10183 16609 10195 16643
rect 11146 16640 11152 16652
rect 10137 16603 10195 16609
rect 10336 16612 11152 16640
rect 10336 16572 10364 16612
rect 10060 16544 10364 16572
rect 10704 16572 10732 16612
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 10873 16575 10931 16581
rect 10873 16572 10885 16575
rect 10704 16544 10885 16572
rect 10873 16541 10885 16544
rect 10919 16541 10931 16575
rect 10873 16535 10931 16541
rect 11241 16575 11299 16581
rect 11241 16541 11253 16575
rect 11287 16572 11299 16575
rect 11348 16572 11376 16680
rect 11606 16668 11612 16720
rect 11664 16708 11670 16720
rect 11664 16680 12388 16708
rect 11664 16668 11670 16680
rect 11514 16600 11520 16652
rect 11572 16600 11578 16652
rect 11287 16544 11376 16572
rect 11532 16572 11560 16600
rect 12360 16581 12388 16680
rect 16592 16649 16620 16748
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 18414 16736 18420 16788
rect 18472 16736 18478 16788
rect 18693 16779 18751 16785
rect 18693 16745 18705 16779
rect 18739 16776 18751 16779
rect 19702 16776 19708 16788
rect 18739 16748 19708 16776
rect 18739 16745 18751 16748
rect 18693 16739 18751 16745
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 25590 16736 25596 16788
rect 25648 16736 25654 16788
rect 18874 16668 18880 16720
rect 18932 16668 18938 16720
rect 25501 16711 25559 16717
rect 25501 16677 25513 16711
rect 25547 16708 25559 16711
rect 25547 16680 26188 16708
rect 25547 16677 25559 16680
rect 25501 16671 25559 16677
rect 26160 16649 26188 16680
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16609 16635 16643
rect 16577 16603 16635 16609
rect 26145 16643 26203 16649
rect 26145 16609 26157 16643
rect 26191 16609 26203 16643
rect 26145 16603 26203 16609
rect 26234 16600 26240 16652
rect 26292 16640 26298 16652
rect 26881 16643 26939 16649
rect 26881 16640 26893 16643
rect 26292 16612 26893 16640
rect 26292 16600 26298 16612
rect 26881 16609 26893 16612
rect 26927 16609 26939 16643
rect 26881 16603 26939 16609
rect 11701 16575 11759 16581
rect 11701 16572 11713 16575
rect 11532 16544 11713 16572
rect 11287 16541 11299 16544
rect 11241 16535 11299 16541
rect 11701 16541 11713 16544
rect 11747 16541 11759 16575
rect 11701 16535 11759 16541
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 11054 16464 11060 16516
rect 11112 16464 11118 16516
rect 11146 16464 11152 16516
rect 11204 16504 11210 16516
rect 11808 16504 11836 16535
rect 12526 16532 12532 16584
rect 12584 16532 12590 16584
rect 16850 16581 16856 16584
rect 16844 16572 16856 16581
rect 16811 16544 16856 16572
rect 16844 16535 16856 16544
rect 16850 16532 16856 16535
rect 16908 16532 16914 16584
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 18141 16575 18199 16581
rect 18141 16572 18153 16575
rect 17368 16544 18153 16572
rect 17368 16532 17374 16544
rect 18141 16541 18153 16544
rect 18187 16541 18199 16575
rect 18141 16535 18199 16541
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16572 18475 16575
rect 19794 16572 19800 16584
rect 18463 16544 19800 16572
rect 18463 16541 18475 16544
rect 18417 16535 18475 16541
rect 11204 16476 11836 16504
rect 18156 16504 18184 16535
rect 19794 16532 19800 16544
rect 19852 16532 19858 16584
rect 25498 16532 25504 16584
rect 25556 16532 25562 16584
rect 25866 16532 25872 16584
rect 25924 16532 25930 16584
rect 18156 16476 18368 16504
rect 11204 16464 11210 16476
rect 5721 16439 5779 16445
rect 5721 16405 5733 16439
rect 5767 16436 5779 16439
rect 5810 16436 5816 16448
rect 5767 16408 5816 16436
rect 5767 16405 5779 16408
rect 5721 16399 5779 16405
rect 5810 16396 5816 16408
rect 5868 16396 5874 16448
rect 6270 16396 6276 16448
rect 6328 16436 6334 16448
rect 7101 16439 7159 16445
rect 7101 16436 7113 16439
rect 6328 16408 7113 16436
rect 6328 16396 6334 16408
rect 7101 16405 7113 16408
rect 7147 16405 7159 16439
rect 7101 16399 7159 16405
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 9677 16439 9735 16445
rect 9677 16436 9689 16439
rect 7708 16408 9689 16436
rect 7708 16396 7714 16408
rect 9677 16405 9689 16408
rect 9723 16405 9735 16439
rect 9677 16399 9735 16405
rect 11425 16439 11483 16445
rect 11425 16405 11437 16439
rect 11471 16436 11483 16439
rect 11514 16436 11520 16448
rect 11471 16408 11520 16436
rect 11471 16405 11483 16408
rect 11425 16399 11483 16405
rect 11514 16396 11520 16408
rect 11572 16396 11578 16448
rect 17957 16439 18015 16445
rect 17957 16405 17969 16439
rect 18003 16436 18015 16439
rect 18230 16436 18236 16448
rect 18003 16408 18236 16436
rect 18003 16405 18015 16408
rect 17957 16399 18015 16405
rect 18230 16396 18236 16408
rect 18288 16396 18294 16448
rect 18340 16436 18368 16476
rect 18506 16464 18512 16516
rect 18564 16464 18570 16516
rect 26789 16507 26847 16513
rect 26789 16473 26801 16507
rect 26835 16504 26847 16507
rect 27126 16507 27184 16513
rect 27126 16504 27138 16507
rect 26835 16476 27138 16504
rect 26835 16473 26847 16476
rect 26789 16467 26847 16473
rect 27126 16473 27138 16476
rect 27172 16473 27184 16507
rect 27126 16467 27184 16473
rect 18709 16439 18767 16445
rect 18709 16436 18721 16439
rect 18340 16408 18721 16436
rect 18709 16405 18721 16408
rect 18755 16405 18767 16439
rect 18709 16399 18767 16405
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 25590 16436 25596 16448
rect 24912 16408 25596 16436
rect 24912 16396 24918 16408
rect 25590 16396 25596 16408
rect 25648 16436 25654 16448
rect 25777 16439 25835 16445
rect 25777 16436 25789 16439
rect 25648 16408 25789 16436
rect 25648 16396 25654 16408
rect 25777 16405 25789 16408
rect 25823 16405 25835 16439
rect 25777 16399 25835 16405
rect 28258 16396 28264 16448
rect 28316 16396 28322 16448
rect 1104 16346 28888 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 28888 16346
rect 1104 16272 28888 16294
rect 5534 16192 5540 16244
rect 5592 16192 5598 16244
rect 6181 16235 6239 16241
rect 6181 16201 6193 16235
rect 6227 16232 6239 16235
rect 7745 16235 7803 16241
rect 6227 16204 6500 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6472 16164 6500 16204
rect 7745 16201 7757 16235
rect 7791 16232 7803 16235
rect 8294 16232 8300 16244
rect 7791 16204 8300 16232
rect 7791 16201 7803 16204
rect 7745 16195 7803 16201
rect 8294 16192 8300 16204
rect 8352 16232 8358 16244
rect 8570 16232 8576 16244
rect 8352 16204 8576 16232
rect 8352 16192 8358 16204
rect 8570 16192 8576 16204
rect 8628 16192 8634 16244
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 10008 16204 10609 16232
rect 10008 16192 10014 16204
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11333 16235 11391 16241
rect 11333 16232 11345 16235
rect 11204 16204 11345 16232
rect 11204 16192 11210 16204
rect 11333 16201 11345 16204
rect 11379 16201 11391 16235
rect 11333 16195 11391 16201
rect 18230 16192 18236 16244
rect 18288 16232 18294 16244
rect 18506 16232 18512 16244
rect 18288 16204 18512 16232
rect 18288 16192 18294 16204
rect 18506 16192 18512 16204
rect 18564 16232 18570 16244
rect 18969 16235 19027 16241
rect 18969 16232 18981 16235
rect 18564 16204 18981 16232
rect 18564 16192 18570 16204
rect 18969 16201 18981 16204
rect 19015 16201 19027 16235
rect 18969 16195 19027 16201
rect 25225 16235 25283 16241
rect 25225 16201 25237 16235
rect 25271 16232 25283 16235
rect 25498 16232 25504 16244
rect 25271 16204 25504 16232
rect 25271 16201 25283 16204
rect 25225 16195 25283 16201
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 28442 16192 28448 16244
rect 28500 16192 28506 16244
rect 6610 16167 6668 16173
rect 6610 16164 6622 16167
rect 4172 16136 6408 16164
rect 6472 16136 6622 16164
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 4172 16105 4200 16136
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 900 16068 1409 16096
rect 900 16056 906 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16065 4215 16099
rect 4413 16099 4471 16105
rect 4413 16096 4425 16099
rect 4157 16059 4215 16065
rect 4264 16068 4425 16096
rect 3418 15988 3424 16040
rect 3476 16028 3482 16040
rect 4264 16028 4292 16068
rect 4413 16065 4425 16068
rect 4459 16065 4471 16099
rect 4413 16059 4471 16065
rect 5810 16056 5816 16108
rect 5868 16056 5874 16108
rect 5994 16056 6000 16108
rect 6052 16056 6058 16108
rect 6380 16105 6408 16136
rect 6610 16133 6622 16136
rect 6656 16133 6668 16167
rect 6610 16127 6668 16133
rect 8205 16167 8263 16173
rect 8205 16133 8217 16167
rect 8251 16164 8263 16167
rect 9490 16164 9496 16176
rect 8251 16136 9496 16164
rect 8251 16133 8263 16136
rect 8205 16127 8263 16133
rect 9490 16124 9496 16136
rect 9548 16124 9554 16176
rect 12158 16124 12164 16176
rect 12216 16164 12222 16176
rect 12314 16167 12372 16173
rect 12314 16164 12326 16167
rect 12216 16136 12326 16164
rect 12216 16124 12222 16136
rect 12314 16133 12326 16136
rect 12360 16133 12372 16167
rect 12314 16127 12372 16133
rect 18138 16124 18144 16176
rect 18196 16164 18202 16176
rect 19153 16167 19211 16173
rect 19153 16164 19165 16167
rect 18196 16136 19165 16164
rect 18196 16124 18202 16136
rect 19153 16133 19165 16136
rect 19199 16164 19211 16167
rect 21450 16164 21456 16176
rect 19199 16136 21456 16164
rect 19199 16133 19211 16136
rect 19153 16127 19211 16133
rect 21450 16124 21456 16136
rect 21508 16124 21514 16176
rect 24029 16167 24087 16173
rect 23676 16136 23980 16164
rect 6365 16099 6423 16105
rect 6365 16065 6377 16099
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 3476 16000 4292 16028
rect 3476 15988 3482 16000
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 3234 15892 3240 15904
rect 1627 15864 3240 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 6380 15892 6408 16059
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 10229 16099 10287 16105
rect 10229 16096 10241 16099
rect 8352 16068 10241 16096
rect 8352 16056 8358 16068
rect 10229 16065 10241 16068
rect 10275 16065 10287 16099
rect 10229 16059 10287 16065
rect 10318 16056 10324 16108
rect 10376 16056 10382 16108
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16096 10471 16099
rect 10594 16096 10600 16108
rect 10459 16068 10600 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 10594 16056 10600 16068
rect 10652 16056 10658 16108
rect 17770 16056 17776 16108
rect 17828 16105 17834 16108
rect 17828 16059 17840 16105
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18322 16096 18328 16108
rect 18095 16068 18328 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 17828 16056 17834 16059
rect 18322 16056 18328 16068
rect 18380 16056 18386 16108
rect 18877 16099 18935 16105
rect 18877 16065 18889 16099
rect 18923 16065 18935 16099
rect 18877 16059 18935 16065
rect 10686 15988 10692 16040
rect 10744 15988 10750 16040
rect 12066 15988 12072 16040
rect 12124 15988 12130 16040
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 18064 16000 18705 16028
rect 8478 15920 8484 15972
rect 8536 15960 8542 15972
rect 10045 15963 10103 15969
rect 10045 15960 10057 15963
rect 8536 15932 10057 15960
rect 8536 15920 8542 15932
rect 10045 15929 10057 15932
rect 10091 15929 10103 15963
rect 10045 15923 10103 15929
rect 7282 15892 7288 15904
rect 6380 15864 7288 15892
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 9030 15852 9036 15904
rect 9088 15892 9094 15904
rect 9493 15895 9551 15901
rect 9493 15892 9505 15895
rect 9088 15864 9505 15892
rect 9088 15852 9094 15864
rect 9493 15861 9505 15864
rect 9539 15861 9551 15895
rect 9493 15855 9551 15861
rect 13449 15895 13507 15901
rect 13449 15861 13461 15895
rect 13495 15892 13507 15895
rect 13722 15892 13728 15904
rect 13495 15864 13728 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 16669 15895 16727 15901
rect 16669 15861 16681 15895
rect 16715 15892 16727 15895
rect 17310 15892 17316 15904
rect 16715 15864 17316 15892
rect 16715 15861 16727 15864
rect 16669 15855 16727 15861
rect 17310 15852 17316 15864
rect 17368 15892 17374 15904
rect 18064 15892 18092 16000
rect 18693 15997 18705 16000
rect 18739 16028 18751 16031
rect 18892 16028 18920 16059
rect 23290 16056 23296 16108
rect 23348 16056 23354 16108
rect 23474 16056 23480 16108
rect 23532 16056 23538 16108
rect 23676 16105 23704 16136
rect 23661 16099 23719 16105
rect 23661 16065 23673 16099
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 23845 16099 23903 16105
rect 23845 16065 23857 16099
rect 23891 16065 23903 16099
rect 23952 16096 23980 16136
rect 24029 16133 24041 16167
rect 24075 16164 24087 16167
rect 24075 16136 24992 16164
rect 24075 16133 24087 16136
rect 24029 16127 24087 16133
rect 24302 16096 24308 16108
rect 23952 16068 24308 16096
rect 23845 16059 23903 16065
rect 18739 16000 18920 16028
rect 18739 15997 18751 16000
rect 18693 15991 18751 15997
rect 22186 15988 22192 16040
rect 22244 16028 22250 16040
rect 23382 16028 23388 16040
rect 22244 16000 23388 16028
rect 22244 15988 22250 16000
rect 23382 15988 23388 16000
rect 23440 16028 23446 16040
rect 23569 16031 23627 16037
rect 23569 16028 23581 16031
rect 23440 16000 23581 16028
rect 23440 15988 23446 16000
rect 23569 15997 23581 16000
rect 23615 15997 23627 16031
rect 23569 15991 23627 15997
rect 23860 15960 23888 16059
rect 24302 16056 24308 16068
rect 24360 16096 24366 16108
rect 24397 16099 24455 16105
rect 24397 16096 24409 16099
rect 24360 16068 24409 16096
rect 24360 16056 24366 16068
rect 24397 16065 24409 16068
rect 24443 16065 24455 16099
rect 24397 16059 24455 16065
rect 24673 16099 24731 16105
rect 24673 16065 24685 16099
rect 24719 16096 24731 16099
rect 24854 16096 24860 16108
rect 24719 16068 24860 16096
rect 24719 16065 24731 16068
rect 24673 16059 24731 16065
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 24964 16105 24992 16136
rect 24949 16099 25007 16105
rect 24949 16065 24961 16099
rect 24995 16065 25007 16099
rect 24949 16059 25007 16065
rect 25041 16099 25099 16105
rect 25041 16065 25053 16099
rect 25087 16065 25099 16099
rect 25041 16059 25099 16065
rect 24213 16031 24271 16037
rect 24213 15997 24225 16031
rect 24259 15997 24271 16031
rect 24213 15991 24271 15997
rect 24581 16031 24639 16037
rect 24581 15997 24593 16031
rect 24627 16028 24639 16031
rect 25056 16028 25084 16059
rect 28258 16056 28264 16108
rect 28316 16056 28322 16108
rect 24627 16000 25084 16028
rect 24627 15997 24639 16000
rect 24581 15991 24639 15997
rect 24228 15960 24256 15991
rect 23860 15932 24256 15960
rect 17368 15864 18092 15892
rect 17368 15852 17374 15864
rect 18138 15852 18144 15904
rect 18196 15852 18202 15904
rect 19150 15852 19156 15904
rect 19208 15852 19214 15904
rect 24228 15892 24256 15932
rect 24765 15963 24823 15969
rect 24765 15929 24777 15963
rect 24811 15960 24823 15963
rect 26510 15960 26516 15972
rect 24811 15932 26516 15960
rect 24811 15929 24823 15932
rect 24765 15923 24823 15929
rect 26510 15920 26516 15932
rect 26568 15920 26574 15972
rect 25222 15892 25228 15904
rect 24228 15864 25228 15892
rect 25222 15852 25228 15864
rect 25280 15852 25286 15904
rect 28166 15852 28172 15904
rect 28224 15852 28230 15904
rect 1104 15802 28888 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 28888 15802
rect 1104 15728 28888 15750
rect 3418 15648 3424 15700
rect 3476 15648 3482 15700
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 7708 15660 8309 15688
rect 7708 15648 7714 15660
rect 8297 15657 8309 15660
rect 8343 15657 8355 15691
rect 8297 15651 8355 15657
rect 11054 15648 11060 15700
rect 11112 15648 11118 15700
rect 11606 15688 11612 15700
rect 11164 15660 11612 15688
rect 8018 15580 8024 15632
rect 8076 15620 8082 15632
rect 11164 15620 11192 15660
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 12621 15691 12679 15697
rect 12621 15688 12633 15691
rect 12584 15660 12633 15688
rect 12584 15648 12590 15660
rect 12621 15657 12633 15660
rect 12667 15657 12679 15691
rect 12621 15651 12679 15657
rect 17681 15691 17739 15697
rect 17681 15657 17693 15691
rect 17727 15688 17739 15691
rect 17770 15688 17776 15700
rect 17727 15660 17776 15688
rect 17727 15657 17739 15660
rect 17681 15651 17739 15657
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 18138 15648 18144 15700
rect 18196 15648 18202 15700
rect 8076 15592 11192 15620
rect 8076 15580 8082 15592
rect 3053 15555 3111 15561
rect 3053 15521 3065 15555
rect 3099 15552 3111 15555
rect 3099 15524 5672 15552
rect 3099 15521 3111 15524
rect 3053 15515 3111 15521
rect 3234 15444 3240 15496
rect 3292 15444 3298 15496
rect 5644 15484 5672 15524
rect 6270 15512 6276 15564
rect 6328 15512 6334 15564
rect 8478 15512 8484 15564
rect 8536 15512 8542 15564
rect 19150 15552 19156 15564
rect 17972 15524 19156 15552
rect 5994 15484 6000 15496
rect 5644 15456 6000 15484
rect 5994 15444 6000 15456
rect 6052 15484 6058 15496
rect 6457 15487 6515 15493
rect 6457 15484 6469 15487
rect 6052 15456 6469 15484
rect 6052 15444 6058 15456
rect 6457 15453 6469 15456
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15484 6791 15487
rect 7282 15484 7288 15496
rect 6779 15456 7288 15484
rect 6779 15453 6791 15456
rect 6733 15447 6791 15453
rect 6472 15348 6500 15447
rect 7282 15444 7288 15456
rect 7340 15484 7346 15496
rect 7340 15456 8524 15484
rect 7340 15444 7346 15456
rect 6641 15419 6699 15425
rect 6641 15385 6653 15419
rect 6687 15416 6699 15419
rect 6978 15419 7036 15425
rect 6978 15416 6990 15419
rect 6687 15388 6990 15416
rect 6687 15385 6699 15388
rect 6641 15379 6699 15385
rect 6978 15385 6990 15388
rect 7024 15385 7036 15419
rect 8294 15416 8300 15428
rect 6978 15379 7036 15385
rect 8128 15388 8300 15416
rect 7834 15348 7840 15360
rect 6472 15320 7840 15348
rect 7834 15308 7840 15320
rect 7892 15348 7898 15360
rect 8018 15348 8024 15360
rect 7892 15320 8024 15348
rect 7892 15308 7898 15320
rect 8018 15308 8024 15320
rect 8076 15308 8082 15360
rect 8128 15357 8156 15388
rect 8294 15376 8300 15388
rect 8352 15376 8358 15428
rect 8496 15416 8524 15456
rect 8570 15444 8576 15496
rect 8628 15444 8634 15496
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15484 10563 15487
rect 10962 15484 10968 15496
rect 10551 15456 10968 15484
rect 10551 15453 10563 15456
rect 10505 15447 10563 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15484 11299 15487
rect 11330 15484 11336 15496
rect 11287 15456 11336 15484
rect 11287 15453 11299 15456
rect 11241 15447 11299 15453
rect 8941 15419 8999 15425
rect 8941 15416 8953 15419
rect 8496 15388 8953 15416
rect 8941 15385 8953 15388
rect 8987 15416 8999 15419
rect 9030 15416 9036 15428
rect 8987 15388 9036 15416
rect 8987 15385 8999 15388
rect 8941 15379 8999 15385
rect 9030 15376 9036 15388
rect 9088 15416 9094 15428
rect 11256 15416 11284 15447
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11514 15493 11520 15496
rect 11508 15447 11520 15493
rect 11514 15444 11520 15447
rect 11572 15444 11578 15496
rect 17972 15493 18000 15524
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15484 17187 15487
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 17175 15456 17785 15484
rect 17175 15453 17187 15456
rect 17129 15447 17187 15453
rect 17773 15453 17785 15456
rect 17819 15453 17831 15487
rect 17773 15447 17831 15453
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15453 18015 15487
rect 17957 15447 18015 15453
rect 18230 15444 18236 15496
rect 18288 15444 18294 15496
rect 19886 15444 19892 15496
rect 19944 15444 19950 15496
rect 19978 15444 19984 15496
rect 20036 15444 20042 15496
rect 20354 15487 20412 15493
rect 20354 15453 20366 15487
rect 20400 15484 20412 15487
rect 20622 15484 20628 15496
rect 20400 15456 20628 15484
rect 20400 15453 20412 15456
rect 20354 15447 20412 15453
rect 9088 15388 11284 15416
rect 9088 15376 9094 15388
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 20165 15419 20223 15425
rect 20165 15416 20177 15419
rect 19392 15388 20177 15416
rect 19392 15376 19398 15388
rect 20165 15385 20177 15388
rect 20211 15385 20223 15419
rect 20165 15379 20223 15385
rect 20254 15376 20260 15428
rect 20312 15376 20318 15428
rect 8113 15351 8171 15357
rect 8113 15317 8125 15351
rect 8159 15317 8171 15351
rect 8113 15311 8171 15317
rect 8757 15351 8815 15357
rect 8757 15317 8769 15351
rect 8803 15348 8815 15351
rect 10502 15348 10508 15360
rect 8803 15320 10508 15348
rect 8803 15317 8815 15320
rect 8757 15311 8815 15317
rect 10502 15308 10508 15320
rect 10560 15308 10566 15360
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 20364 15348 20392 15447
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 20806 15444 20812 15496
rect 20864 15484 20870 15496
rect 21453 15487 21511 15493
rect 21453 15484 21465 15487
rect 20864 15456 21465 15484
rect 20864 15444 20870 15456
rect 21453 15453 21465 15456
rect 21499 15453 21511 15487
rect 21453 15447 21511 15453
rect 21542 15444 21548 15496
rect 21600 15484 21606 15496
rect 21600 15456 21645 15484
rect 21600 15444 21606 15456
rect 19484 15320 20392 15348
rect 20533 15351 20591 15357
rect 19484 15308 19490 15320
rect 20533 15317 20545 15351
rect 20579 15348 20591 15351
rect 21726 15348 21732 15360
rect 20579 15320 21732 15348
rect 20579 15317 20591 15320
rect 20533 15311 20591 15317
rect 21726 15308 21732 15320
rect 21784 15308 21790 15360
rect 21821 15351 21879 15357
rect 21821 15317 21833 15351
rect 21867 15348 21879 15351
rect 22094 15348 22100 15360
rect 21867 15320 22100 15348
rect 21867 15317 21879 15320
rect 21821 15311 21879 15317
rect 22094 15308 22100 15320
rect 22152 15308 22158 15360
rect 1104 15258 28888 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 28888 15258
rect 1104 15184 28888 15206
rect 8478 15104 8484 15156
rect 8536 15144 8542 15156
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 8536 15116 8677 15144
rect 8536 15104 8542 15116
rect 8665 15113 8677 15116
rect 8711 15113 8723 15147
rect 8665 15107 8723 15113
rect 10413 15147 10471 15153
rect 10413 15113 10425 15147
rect 10459 15144 10471 15147
rect 10686 15144 10692 15156
rect 10459 15116 10692 15144
rect 10459 15113 10471 15116
rect 10413 15107 10471 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 10962 15104 10968 15156
rect 11020 15104 11026 15156
rect 22465 15147 22523 15153
rect 14108 15116 14780 15144
rect 7300 15048 9076 15076
rect 7300 15017 7328 15048
rect 7558 15017 7564 15020
rect 7285 15011 7343 15017
rect 7285 14977 7297 15011
rect 7331 14977 7343 15011
rect 7285 14971 7343 14977
rect 7552 14971 7564 15017
rect 7558 14968 7564 14971
rect 7616 14968 7622 15020
rect 9048 14952 9076 15048
rect 10502 15036 10508 15088
rect 10560 15036 10566 15088
rect 13722 15036 13728 15088
rect 13780 15076 13786 15088
rect 14108 15085 14136 15116
rect 14093 15079 14151 15085
rect 14093 15076 14105 15079
rect 13780 15048 14105 15076
rect 13780 15036 13786 15048
rect 14093 15045 14105 15048
rect 14139 15045 14151 15079
rect 14093 15039 14151 15045
rect 14277 15079 14335 15085
rect 14277 15045 14289 15079
rect 14323 15076 14335 15079
rect 14553 15079 14611 15085
rect 14553 15076 14565 15079
rect 14323 15048 14565 15076
rect 14323 15045 14335 15048
rect 14277 15039 14335 15045
rect 14553 15045 14565 15048
rect 14599 15045 14611 15079
rect 14553 15039 14611 15045
rect 9300 15011 9358 15017
rect 9300 14977 9312 15011
rect 9346 15008 9358 15011
rect 9674 15008 9680 15020
rect 9346 14980 9680 15008
rect 9346 14977 9358 14980
rect 9300 14971 9358 14977
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 10778 14968 10784 15020
rect 10836 14968 10842 15020
rect 12526 14968 12532 15020
rect 12584 15008 12590 15020
rect 13446 15008 13452 15020
rect 12584 14980 13452 15008
rect 12584 14968 12590 14980
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 13630 14968 13636 15020
rect 13688 15008 13694 15020
rect 14752 15017 14780 15116
rect 22465 15113 22477 15147
rect 22511 15144 22523 15147
rect 23290 15144 23296 15156
rect 22511 15116 23296 15144
rect 22511 15113 22523 15116
rect 22465 15107 22523 15113
rect 23290 15104 23296 15116
rect 23348 15104 23354 15156
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 17681 15079 17739 15085
rect 17681 15076 17693 15079
rect 17276 15048 17693 15076
rect 17276 15036 17282 15048
rect 17681 15045 17693 15048
rect 17727 15045 17739 15079
rect 17681 15039 17739 15045
rect 22094 15036 22100 15088
rect 22152 15036 22158 15088
rect 22186 15036 22192 15088
rect 22244 15036 22250 15088
rect 13909 15011 13967 15017
rect 13909 15008 13921 15011
rect 13688 14980 13921 15008
rect 13688 14968 13694 14980
rect 13909 14977 13921 14980
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 14369 15011 14427 15017
rect 14369 14977 14381 15011
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 14737 15011 14795 15017
rect 14737 14977 14749 15011
rect 14783 14977 14795 15011
rect 14737 14971 14795 14977
rect 9030 14900 9036 14952
rect 9088 14900 9094 14952
rect 10594 14900 10600 14952
rect 10652 14900 10658 14952
rect 13538 14900 13544 14952
rect 13596 14900 13602 14952
rect 13817 14875 13875 14881
rect 13817 14841 13829 14875
rect 13863 14872 13875 14875
rect 14384 14872 14412 14971
rect 14660 14940 14688 14971
rect 14918 14968 14924 15020
rect 14976 14968 14982 15020
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 17497 15011 17555 15017
rect 17497 15008 17509 15011
rect 17368 14980 17509 15008
rect 17368 14968 17374 14980
rect 17497 14977 17509 14980
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 21726 14968 21732 15020
rect 21784 15008 21790 15020
rect 21913 15011 21971 15017
rect 21913 15008 21925 15011
rect 21784 14980 21925 15008
rect 21784 14968 21790 14980
rect 21913 14977 21925 14980
rect 21959 14977 21971 15011
rect 21913 14971 21971 14977
rect 22281 15011 22339 15017
rect 22281 14977 22293 15011
rect 22327 15008 22339 15011
rect 23474 15008 23480 15020
rect 22327 14980 23480 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 23474 14968 23480 14980
rect 23532 14968 23538 15020
rect 14829 14943 14887 14949
rect 14829 14940 14841 14943
rect 14660 14912 14841 14940
rect 14829 14909 14841 14912
rect 14875 14909 14887 14943
rect 14829 14903 14887 14909
rect 13863 14844 14412 14872
rect 13863 14841 13875 14844
rect 13817 14835 13875 14841
rect 10318 14764 10324 14816
rect 10376 14804 10382 14816
rect 10505 14807 10563 14813
rect 10505 14804 10517 14807
rect 10376 14776 10517 14804
rect 10376 14764 10382 14776
rect 10505 14773 10517 14776
rect 10551 14773 10563 14807
rect 10505 14767 10563 14773
rect 14369 14807 14427 14813
rect 14369 14773 14381 14807
rect 14415 14804 14427 14807
rect 16206 14804 16212 14816
rect 14415 14776 16212 14804
rect 14415 14773 14427 14776
rect 14369 14767 14427 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 17865 14807 17923 14813
rect 17865 14773 17877 14807
rect 17911 14804 17923 14807
rect 18322 14804 18328 14816
rect 17911 14776 18328 14804
rect 17911 14773 17923 14776
rect 17865 14767 17923 14773
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 1104 14714 28888 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 28888 14714
rect 1104 14640 28888 14662
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7616 14572 7665 14600
rect 7616 14560 7622 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 7653 14563 7711 14569
rect 9674 14560 9680 14612
rect 9732 14560 9738 14612
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 13780 14572 14197 14600
rect 13780 14560 13786 14572
rect 14185 14569 14197 14572
rect 14231 14569 14243 14603
rect 14185 14563 14243 14569
rect 18877 14603 18935 14609
rect 18877 14569 18889 14603
rect 18923 14600 18935 14603
rect 19334 14600 19340 14612
rect 18923 14572 19340 14600
rect 18923 14569 18935 14572
rect 18877 14563 18935 14569
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 19797 14603 19855 14609
rect 19797 14569 19809 14603
rect 19843 14600 19855 14603
rect 19978 14600 19984 14612
rect 19843 14572 19984 14600
rect 19843 14569 19855 14572
rect 19797 14563 19855 14569
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 13354 14492 13360 14544
rect 13412 14532 13418 14544
rect 13630 14532 13636 14544
rect 13412 14504 13636 14532
rect 13412 14492 13418 14504
rect 13630 14492 13636 14504
rect 13688 14532 13694 14544
rect 14918 14532 14924 14544
rect 13688 14504 14924 14532
rect 13688 14492 13694 14504
rect 8478 14424 8484 14476
rect 8536 14464 8542 14476
rect 8941 14467 8999 14473
rect 8941 14464 8953 14467
rect 8536 14436 8953 14464
rect 8536 14424 8542 14436
rect 8941 14433 8953 14436
rect 8987 14433 8999 14467
rect 8941 14427 8999 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 9631 14436 10057 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 10045 14433 10057 14436
rect 10091 14433 10103 14467
rect 10045 14427 10103 14433
rect 13464 14436 13676 14464
rect 13464 14408 13492 14436
rect 7834 14356 7840 14408
rect 7892 14356 7898 14408
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14396 8079 14399
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 8067 14368 8125 14396
rect 8067 14365 8079 14368
rect 8021 14359 8079 14365
rect 8113 14365 8125 14368
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8665 14399 8723 14405
rect 8665 14396 8677 14399
rect 8352 14368 8677 14396
rect 8352 14356 8358 14368
rect 8665 14365 8677 14368
rect 8711 14365 8723 14399
rect 8665 14359 8723 14365
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 9824 14368 9873 14396
rect 9824 14356 9830 14368
rect 9861 14365 9873 14368
rect 9907 14396 9919 14399
rect 10226 14396 10232 14408
rect 9907 14368 10232 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 13446 14356 13452 14408
rect 13504 14356 13510 14408
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14365 13599 14399
rect 13648 14396 13676 14436
rect 14384 14405 14412 14504
rect 14918 14492 14924 14504
rect 14976 14492 14982 14544
rect 19702 14532 19708 14544
rect 18708 14504 19708 14532
rect 18230 14464 18236 14476
rect 17052 14436 18236 14464
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13648 14368 14105 14396
rect 13541 14359 13599 14365
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14365 14427 14399
rect 14369 14359 14427 14365
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 13354 14288 13360 14340
rect 13412 14328 13418 14340
rect 13556 14328 13584 14359
rect 13412 14300 13584 14328
rect 13412 14288 13418 14300
rect 13630 14288 13636 14340
rect 13688 14288 13694 14340
rect 13725 14331 13783 14337
rect 13725 14297 13737 14331
rect 13771 14328 13783 14331
rect 14568 14328 14596 14359
rect 16942 14356 16948 14408
rect 17000 14356 17006 14408
rect 17052 14405 17080 14436
rect 18230 14424 18236 14436
rect 18288 14424 18294 14476
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 17218 14356 17224 14408
rect 17276 14356 17282 14408
rect 17310 14356 17316 14408
rect 17368 14356 17374 14408
rect 18322 14356 18328 14408
rect 18380 14356 18386 14408
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 18708 14405 18736 14504
rect 19702 14492 19708 14504
rect 19760 14492 19766 14544
rect 19886 14492 19892 14544
rect 19944 14532 19950 14544
rect 20625 14535 20683 14541
rect 20625 14532 20637 14535
rect 19944 14504 20637 14532
rect 19944 14492 19950 14504
rect 20625 14501 20637 14504
rect 20671 14501 20683 14535
rect 20625 14495 20683 14501
rect 20806 14492 20812 14544
rect 20864 14492 20870 14544
rect 19334 14424 19340 14476
rect 19392 14424 19398 14476
rect 20254 14464 20260 14476
rect 19444 14436 20260 14464
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18472 14368 18613 14396
rect 18472 14356 18478 14368
rect 18601 14365 18613 14368
rect 18647 14365 18659 14399
rect 18601 14359 18659 14365
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 15470 14328 15476 14340
rect 13771 14300 14596 14328
rect 14660 14300 15476 14328
rect 13771 14297 13783 14300
rect 13725 14291 13783 14297
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 13740 14260 13768 14291
rect 13504 14232 13768 14260
rect 13909 14263 13967 14269
rect 13504 14220 13510 14232
rect 13909 14229 13921 14263
rect 13955 14260 13967 14263
rect 14660 14260 14688 14300
rect 15470 14288 15476 14300
rect 15528 14288 15534 14340
rect 17497 14331 17555 14337
rect 17497 14297 17509 14331
rect 17543 14328 17555 14331
rect 18509 14331 18567 14337
rect 18509 14328 18521 14331
rect 17543 14300 18521 14328
rect 17543 14297 17555 14300
rect 17497 14291 17555 14297
rect 18509 14297 18521 14300
rect 18555 14297 18567 14331
rect 18616 14328 18644 14359
rect 18874 14356 18880 14408
rect 18932 14396 18938 14408
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 18932 14368 19257 14396
rect 18932 14356 18938 14368
rect 19245 14365 19257 14368
rect 19291 14396 19303 14399
rect 19444 14396 19472 14436
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 19291 14368 19472 14396
rect 19521 14399 19579 14405
rect 19291 14365 19303 14368
rect 19245 14359 19303 14365
rect 19521 14365 19533 14399
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14396 19671 14399
rect 19702 14396 19708 14408
rect 19659 14368 19708 14396
rect 19659 14365 19671 14368
rect 19613 14359 19671 14365
rect 19536 14328 19564 14359
rect 19702 14356 19708 14368
rect 19760 14356 19766 14408
rect 18616 14300 19564 14328
rect 21085 14331 21143 14337
rect 18509 14291 18567 14297
rect 21085 14297 21097 14331
rect 21131 14328 21143 14331
rect 21542 14328 21548 14340
rect 21131 14300 21548 14328
rect 21131 14297 21143 14300
rect 21085 14291 21143 14297
rect 21542 14288 21548 14300
rect 21600 14288 21606 14340
rect 13955 14232 14688 14260
rect 14737 14263 14795 14269
rect 13955 14229 13967 14232
rect 13909 14223 13967 14229
rect 14737 14229 14749 14263
rect 14783 14260 14795 14263
rect 15286 14260 15292 14272
rect 14783 14232 15292 14260
rect 14783 14229 14795 14232
rect 14737 14223 14795 14229
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 1104 14170 28888 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 28888 14170
rect 1104 14096 28888 14118
rect 25590 14016 25596 14068
rect 25648 14016 25654 14068
rect 18690 13948 18696 14000
rect 18748 13948 18754 14000
rect 16206 13880 16212 13932
rect 16264 13920 16270 13932
rect 25133 13923 25191 13929
rect 25133 13920 25145 13923
rect 16264 13892 25145 13920
rect 16264 13880 16270 13892
rect 25133 13889 25145 13892
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 25314 13880 25320 13932
rect 25372 13880 25378 13932
rect 25682 13880 25688 13932
rect 25740 13880 25746 13932
rect 24949 13855 25007 13861
rect 24949 13821 24961 13855
rect 24995 13852 25007 13855
rect 25406 13852 25412 13864
rect 24995 13824 25412 13852
rect 24995 13821 25007 13824
rect 24949 13815 25007 13821
rect 25406 13812 25412 13824
rect 25464 13812 25470 13864
rect 17218 13676 17224 13728
rect 17276 13676 17282 13728
rect 24854 13676 24860 13728
rect 24912 13676 24918 13728
rect 25038 13676 25044 13728
rect 25096 13676 25102 13728
rect 1104 13626 28888 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 28888 13626
rect 1104 13552 28888 13574
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 13412 13484 13737 13512
rect 13412 13472 13418 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15528 13484 16313 13512
rect 15528 13472 15534 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 24489 13515 24547 13521
rect 24489 13481 24501 13515
rect 24535 13512 24547 13515
rect 25038 13512 25044 13524
rect 24535 13484 25044 13512
rect 24535 13481 24547 13484
rect 24489 13475 24547 13481
rect 25038 13472 25044 13484
rect 25096 13472 25102 13524
rect 25682 13472 25688 13524
rect 25740 13512 25746 13524
rect 26145 13515 26203 13521
rect 26145 13512 26157 13515
rect 25740 13484 26157 13512
rect 25740 13472 25746 13484
rect 26145 13481 26157 13484
rect 26191 13512 26203 13515
rect 26191 13484 26832 13512
rect 26191 13481 26203 13484
rect 26145 13475 26203 13481
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 12345 13379 12403 13385
rect 12345 13376 12357 13379
rect 12124 13348 12357 13376
rect 12124 13336 12130 13348
rect 12345 13345 12357 13348
rect 12391 13345 12403 13379
rect 12345 13339 12403 13345
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13376 15439 13379
rect 16758 13376 16764 13388
rect 15427 13348 16764 13376
rect 15427 13345 15439 13348
rect 15381 13339 15439 13345
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 21818 13376 21824 13388
rect 17236 13348 21824 13376
rect 17236 13320 17264 13348
rect 21818 13336 21824 13348
rect 21876 13376 21882 13388
rect 26804 13385 26832 13484
rect 24765 13379 24823 13385
rect 24765 13376 24777 13379
rect 21876 13348 24777 13376
rect 21876 13336 21882 13348
rect 24765 13345 24777 13348
rect 24811 13345 24823 13379
rect 24765 13339 24823 13345
rect 26789 13379 26847 13385
rect 26789 13345 26801 13379
rect 26835 13345 26847 13379
rect 26789 13339 26847 13345
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 15470 13268 15476 13320
rect 15528 13268 15534 13320
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13308 15899 13311
rect 17129 13311 17187 13317
rect 15887 13280 16528 13308
rect 15887 13277 15899 13280
rect 15841 13271 15899 13277
rect 12618 13249 12624 13252
rect 12612 13203 12624 13249
rect 12618 13200 12624 13203
rect 12676 13200 12682 13252
rect 15304 13240 15332 13268
rect 15580 13240 15608 13271
rect 16500 13249 16528 13280
rect 17129 13277 17141 13311
rect 17175 13308 17187 13311
rect 17218 13308 17224 13320
rect 17175 13280 17224 13308
rect 17175 13277 17187 13280
rect 17129 13271 17187 13277
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 21450 13308 21456 13320
rect 20772 13280 21456 13308
rect 20772 13268 20778 13280
rect 21450 13268 21456 13280
rect 21508 13308 21514 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 21508 13280 21557 13308
rect 21508 13268 21514 13280
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 21545 13271 21603 13277
rect 21726 13268 21732 13320
rect 21784 13268 21790 13320
rect 24486 13268 24492 13320
rect 24544 13268 24550 13320
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13277 24731 13311
rect 24673 13271 24731 13277
rect 16269 13243 16327 13249
rect 16269 13240 16281 13243
rect 15304 13212 16281 13240
rect 16269 13209 16281 13212
rect 16315 13209 16327 13243
rect 16269 13203 16327 13209
rect 16485 13243 16543 13249
rect 16485 13209 16497 13243
rect 16531 13240 16543 13243
rect 16574 13240 16580 13252
rect 16531 13212 16580 13240
rect 16531 13209 16543 13212
rect 16485 13203 16543 13209
rect 16574 13200 16580 13212
rect 16632 13240 16638 13252
rect 17034 13240 17040 13252
rect 16632 13212 17040 13240
rect 16632 13200 16638 13212
rect 17034 13200 17040 13212
rect 17092 13200 17098 13252
rect 24688 13240 24716 13271
rect 24854 13268 24860 13320
rect 24912 13308 24918 13320
rect 25021 13311 25079 13317
rect 25021 13308 25033 13311
rect 24912 13280 25033 13308
rect 24912 13268 24918 13280
rect 25021 13277 25033 13280
rect 25067 13277 25079 13311
rect 25021 13271 25079 13277
rect 26237 13243 26295 13249
rect 26237 13240 26249 13243
rect 24688 13212 26249 13240
rect 26237 13209 26249 13212
rect 26283 13209 26295 13243
rect 26237 13203 26295 13209
rect 15470 13132 15476 13184
rect 15528 13172 15534 13184
rect 15657 13175 15715 13181
rect 15657 13172 15669 13175
rect 15528 13144 15669 13172
rect 15528 13132 15534 13144
rect 15657 13141 15669 13144
rect 15703 13141 15715 13175
rect 15657 13135 15715 13141
rect 16022 13132 16028 13184
rect 16080 13132 16086 13184
rect 16114 13132 16120 13184
rect 16172 13132 16178 13184
rect 21637 13175 21695 13181
rect 21637 13141 21649 13175
rect 21683 13172 21695 13175
rect 22002 13172 22008 13184
rect 21683 13144 22008 13172
rect 21683 13141 21695 13144
rect 21637 13135 21695 13141
rect 22002 13132 22008 13144
rect 22060 13132 22066 13184
rect 1104 13082 28888 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 28888 13082
rect 1104 13008 28888 13030
rect 23201 12971 23259 12977
rect 23201 12937 23213 12971
rect 23247 12937 23259 12971
rect 23201 12931 23259 12937
rect 16022 12860 16028 12912
rect 16080 12900 16086 12912
rect 16669 12903 16727 12909
rect 16669 12900 16681 12903
rect 16080 12872 16681 12900
rect 16080 12860 16086 12872
rect 16669 12869 16681 12872
rect 16715 12869 16727 12903
rect 16669 12863 16727 12869
rect 21284 12872 21956 12900
rect 16114 12792 16120 12844
rect 16172 12832 16178 12844
rect 21284 12841 21312 12872
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 16172 12804 17049 12832
rect 16172 12792 16178 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 21269 12835 21327 12841
rect 21269 12801 21281 12835
rect 21315 12801 21327 12835
rect 21269 12795 21327 12801
rect 21818 12792 21824 12844
rect 21876 12792 21882 12844
rect 21928 12832 21956 12872
rect 22002 12860 22008 12912
rect 22060 12909 22066 12912
rect 22060 12903 22124 12909
rect 22060 12869 22078 12903
rect 22112 12869 22124 12903
rect 22060 12863 22124 12869
rect 22060 12860 22066 12863
rect 22370 12832 22376 12844
rect 21928 12804 22376 12832
rect 22370 12792 22376 12804
rect 22428 12792 22434 12844
rect 23216 12832 23244 12931
rect 23382 12928 23388 12980
rect 23440 12928 23446 12980
rect 25225 12971 25283 12977
rect 25225 12937 25237 12971
rect 25271 12968 25283 12971
rect 25314 12968 25320 12980
rect 25271 12940 25320 12968
rect 25271 12937 25283 12940
rect 25225 12931 25283 12937
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 25590 12928 25596 12980
rect 25648 12928 25654 12980
rect 25608 12900 25636 12928
rect 24780 12872 25636 12900
rect 23290 12832 23296 12844
rect 23216 12804 23296 12832
rect 23290 12792 23296 12804
rect 23348 12792 23354 12844
rect 24780 12841 24808 12872
rect 24765 12835 24823 12841
rect 24765 12801 24777 12835
rect 24811 12801 24823 12835
rect 24765 12795 24823 12801
rect 25590 12792 25596 12844
rect 25648 12792 25654 12844
rect 16942 12724 16948 12776
rect 17000 12724 17006 12776
rect 21358 12724 21364 12776
rect 21416 12724 21422 12776
rect 24673 12767 24731 12773
rect 24673 12733 24685 12767
rect 24719 12764 24731 12767
rect 24854 12764 24860 12776
rect 24719 12736 24860 12764
rect 24719 12733 24731 12736
rect 24673 12727 24731 12733
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 25501 12767 25559 12773
rect 25501 12764 25513 12767
rect 25148 12736 25513 12764
rect 17037 12699 17095 12705
rect 17037 12665 17049 12699
rect 17083 12696 17095 12699
rect 17954 12696 17960 12708
rect 17083 12668 17960 12696
rect 17083 12665 17095 12668
rect 17037 12659 17095 12665
rect 17954 12656 17960 12668
rect 18012 12656 18018 12708
rect 21634 12656 21640 12708
rect 21692 12656 21698 12708
rect 25148 12705 25176 12736
rect 25501 12733 25513 12736
rect 25547 12733 25559 12767
rect 25501 12727 25559 12733
rect 25133 12699 25191 12705
rect 25133 12665 25145 12699
rect 25179 12665 25191 12699
rect 25133 12659 25191 12665
rect 1104 12538 28888 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 28888 12538
rect 1104 12464 28888 12486
rect 11514 12384 11520 12436
rect 11572 12424 11578 12436
rect 12618 12424 12624 12436
rect 11572 12396 12624 12424
rect 11572 12384 11578 12396
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 16942 12424 16948 12436
rect 16347 12396 16948 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 21726 12384 21732 12436
rect 21784 12424 21790 12436
rect 22005 12427 22063 12433
rect 22005 12424 22017 12427
rect 21784 12396 22017 12424
rect 21784 12384 21790 12396
rect 22005 12393 22017 12396
rect 22051 12393 22063 12427
rect 22005 12387 22063 12393
rect 22370 12384 22376 12436
rect 22428 12424 22434 12436
rect 23382 12424 23388 12436
rect 22428 12396 23388 12424
rect 22428 12384 22434 12396
rect 23382 12384 23388 12396
rect 23440 12384 23446 12436
rect 21542 12316 21548 12368
rect 21600 12356 21606 12368
rect 23201 12359 23259 12365
rect 23201 12356 23213 12359
rect 21600 12328 23213 12356
rect 21600 12316 21606 12328
rect 23201 12325 23213 12328
rect 23247 12325 23259 12359
rect 23201 12319 23259 12325
rect 9784 12260 12434 12288
rect 9784 12232 9812 12260
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12220 10011 12223
rect 11698 12220 11704 12232
rect 9999 12192 11704 12220
rect 9999 12189 10011 12192
rect 9953 12183 10011 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 12406 12220 12434 12260
rect 21450 12248 21456 12300
rect 21508 12248 21514 12300
rect 22649 12291 22707 12297
rect 22649 12257 22661 12291
rect 22695 12288 22707 12291
rect 22695 12260 23244 12288
rect 22695 12257 22707 12260
rect 22649 12251 22707 12257
rect 12805 12223 12863 12229
rect 12805 12220 12817 12223
rect 12406 12192 12817 12220
rect 12805 12189 12817 12192
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 13446 12220 13452 12232
rect 13035 12192 13452 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 16209 12223 16267 12229
rect 16209 12220 16221 12223
rect 15252 12192 16221 12220
rect 15252 12180 15258 12192
rect 16209 12189 16221 12192
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 21545 12223 21603 12229
rect 21545 12189 21557 12223
rect 21591 12220 21603 12223
rect 21634 12220 21640 12232
rect 21591 12192 21640 12220
rect 21591 12189 21603 12192
rect 21545 12183 21603 12189
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 22278 12180 22284 12232
rect 22336 12220 22342 12232
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 22336 12192 22845 12220
rect 22336 12180 22342 12192
rect 22833 12189 22845 12192
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 23014 12180 23020 12232
rect 23072 12180 23078 12232
rect 23216 12220 23244 12260
rect 23290 12248 23296 12300
rect 23348 12248 23354 12300
rect 24486 12220 24492 12232
rect 23216 12192 24492 12220
rect 24486 12180 24492 12192
rect 24544 12180 24550 12232
rect 22465 12155 22523 12161
rect 22465 12152 22477 12155
rect 21928 12124 22477 12152
rect 9582 12044 9588 12096
rect 9640 12044 9646 12096
rect 21928 12093 21956 12124
rect 22465 12121 22477 12124
rect 22511 12121 22523 12155
rect 22465 12115 22523 12121
rect 21913 12087 21971 12093
rect 21913 12053 21925 12087
rect 21959 12053 21971 12087
rect 21913 12047 21971 12053
rect 22370 12044 22376 12096
rect 22428 12044 22434 12096
rect 1104 11994 28888 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 28888 11994
rect 1104 11920 28888 11942
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 16574 11880 16580 11892
rect 15703 11852 16580 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 9392 11815 9450 11821
rect 9392 11781 9404 11815
rect 9438 11812 9450 11815
rect 9582 11812 9588 11824
rect 9438 11784 9588 11812
rect 9438 11781 9450 11784
rect 9392 11775 9450 11781
rect 9582 11772 9588 11784
rect 9640 11772 9646 11824
rect 16114 11812 16120 11824
rect 15304 11784 16120 11812
rect 15304 11753 15332 11784
rect 16114 11772 16120 11784
rect 16172 11772 16178 11824
rect 16206 11772 16212 11824
rect 16264 11772 16270 11824
rect 16758 11772 16764 11824
rect 16816 11812 16822 11824
rect 21174 11812 21180 11824
rect 16816 11784 21180 11812
rect 16816 11772 16822 11784
rect 21174 11772 21180 11784
rect 21232 11812 21238 11824
rect 23014 11812 23020 11824
rect 21232 11784 23020 11812
rect 21232 11772 21238 11784
rect 23014 11772 23020 11784
rect 23072 11772 23078 11824
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15746 11704 15752 11756
rect 15804 11704 15810 11756
rect 18414 11704 18420 11756
rect 18472 11704 18478 11756
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 9088 11648 9137 11676
rect 9088 11636 9094 11648
rect 9125 11645 9137 11648
rect 9171 11645 9183 11679
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 9125 11639 9183 11645
rect 10520 11648 12081 11676
rect 10520 11552 10548 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 17037 11679 17095 11685
rect 17037 11676 17049 11679
rect 16540 11648 17049 11676
rect 16540 11636 16546 11648
rect 17037 11645 17049 11648
rect 17083 11676 17095 11679
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 17083 11648 18521 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 18509 11645 18521 11648
rect 18555 11676 18567 11679
rect 18782 11676 18788 11688
rect 18555 11648 18788 11676
rect 18555 11645 18567 11648
rect 18509 11639 18567 11645
rect 18782 11636 18788 11648
rect 18840 11636 18846 11688
rect 16022 11568 16028 11620
rect 16080 11568 16086 11620
rect 18046 11568 18052 11620
rect 18104 11568 18110 11620
rect 10502 11500 10508 11552
rect 10560 11500 10566 11552
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 11517 11543 11575 11549
rect 11517 11540 11529 11543
rect 11388 11512 11529 11540
rect 11388 11500 11394 11512
rect 11517 11509 11529 11512
rect 11563 11509 11575 11543
rect 11517 11503 11575 11509
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 15289 11543 15347 11549
rect 15289 11540 15301 11543
rect 15160 11512 15301 11540
rect 15160 11500 15166 11512
rect 15289 11509 15301 11512
rect 15335 11509 15347 11543
rect 15289 11503 15347 11509
rect 1104 11450 28888 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 28888 11450
rect 1104 11376 28888 11398
rect 11698 11296 11704 11348
rect 11756 11296 11762 11348
rect 13446 11296 13452 11348
rect 13504 11296 13510 11348
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 15528 11308 16313 11336
rect 15528 11296 15534 11308
rect 16301 11305 16313 11308
rect 16347 11305 16359 11339
rect 16301 11299 16359 11305
rect 21450 11296 21456 11348
rect 21508 11336 21514 11348
rect 21545 11339 21603 11345
rect 21545 11336 21557 11339
rect 21508 11308 21557 11336
rect 21508 11296 21514 11308
rect 21545 11305 21557 11308
rect 21591 11305 21603 11339
rect 21545 11299 21603 11305
rect 10321 11271 10379 11277
rect 10321 11237 10333 11271
rect 10367 11268 10379 11271
rect 15381 11271 15439 11277
rect 10367 11240 11100 11268
rect 10367 11237 10379 11240
rect 10321 11231 10379 11237
rect 11072 11209 11100 11240
rect 15381 11237 15393 11271
rect 15427 11268 15439 11271
rect 16574 11268 16580 11280
rect 15427 11240 15976 11268
rect 15427 11237 15439 11240
rect 15381 11231 15439 11237
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 12066 11160 12072 11212
rect 12124 11160 12130 11212
rect 15102 11160 15108 11212
rect 15160 11160 15166 11212
rect 15948 11209 15976 11240
rect 16132 11240 16580 11268
rect 15933 11203 15991 11209
rect 15933 11169 15945 11203
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 16022 11160 16028 11212
rect 16080 11160 16086 11212
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11132 8999 11135
rect 9030 11132 9036 11144
rect 8987 11104 9036 11132
rect 8987 11101 8999 11104
rect 8941 11095 8999 11101
rect 9030 11092 9036 11104
rect 9088 11132 9094 11144
rect 15013 11135 15071 11141
rect 9088 11104 9352 11132
rect 9088 11092 9094 11104
rect 9324 11076 9352 11104
rect 15013 11101 15025 11135
rect 15059 11132 15071 11135
rect 15194 11132 15200 11144
rect 15059 11104 15200 11132
rect 15059 11101 15071 11104
rect 15013 11095 15071 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11132 15899 11135
rect 16132 11132 16160 11240
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 21634 11228 21640 11280
rect 21692 11268 21698 11280
rect 21692 11240 22600 11268
rect 21692 11228 21698 11240
rect 21266 11160 21272 11212
rect 21324 11200 21330 11212
rect 21910 11200 21916 11212
rect 21324 11172 21916 11200
rect 21324 11160 21330 11172
rect 15887 11104 16160 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 16482 11092 16488 11144
rect 16540 11092 16546 11144
rect 16577 11135 16635 11141
rect 16577 11101 16589 11135
rect 16623 11101 16635 11135
rect 16577 11095 16635 11101
rect 9214 11073 9220 11076
rect 9208 11027 9220 11073
rect 9214 11024 9220 11027
rect 9272 11024 9278 11076
rect 9306 11024 9312 11076
rect 9364 11024 9370 11076
rect 12336 11067 12394 11073
rect 12336 11033 12348 11067
rect 12382 11064 12394 11067
rect 12894 11064 12900 11076
rect 12382 11036 12900 11064
rect 12382 11033 12394 11036
rect 12336 11027 12394 11033
rect 12894 11024 12900 11036
rect 12952 11024 12958 11076
rect 15746 11024 15752 11076
rect 15804 11064 15810 11076
rect 16592 11064 16620 11095
rect 21358 11092 21364 11144
rect 21416 11132 21422 11144
rect 21729 11135 21787 11141
rect 21729 11132 21741 11135
rect 21416 11104 21741 11132
rect 21416 11092 21422 11104
rect 21729 11101 21741 11104
rect 21775 11101 21787 11135
rect 21836 11132 21864 11172
rect 21910 11160 21916 11172
rect 21968 11160 21974 11212
rect 22572 11209 22600 11240
rect 22465 11203 22523 11209
rect 22465 11200 22477 11203
rect 22112 11172 22477 11200
rect 22112 11141 22140 11172
rect 22465 11169 22477 11172
rect 22511 11169 22523 11203
rect 22465 11163 22523 11169
rect 22557 11203 22615 11209
rect 22557 11169 22569 11203
rect 22603 11169 22615 11203
rect 22557 11163 22615 11169
rect 22741 11203 22799 11209
rect 22741 11169 22753 11203
rect 22787 11200 22799 11203
rect 24486 11200 24492 11212
rect 22787 11172 24492 11200
rect 22787 11169 22799 11172
rect 22741 11163 22799 11169
rect 24486 11160 24492 11172
rect 24544 11160 24550 11212
rect 22097 11135 22155 11141
rect 22097 11132 22109 11135
rect 21836 11104 22109 11132
rect 21729 11095 21787 11101
rect 22097 11101 22109 11104
rect 22143 11101 22155 11135
rect 22097 11095 22155 11101
rect 22278 11092 22284 11144
rect 22336 11092 22342 11144
rect 22373 11135 22431 11141
rect 22373 11101 22385 11135
rect 22419 11101 22431 11135
rect 22373 11095 22431 11101
rect 15804 11036 16620 11064
rect 15804 11024 15810 11036
rect 21542 11024 21548 11076
rect 21600 11064 21606 11076
rect 21821 11067 21879 11073
rect 21821 11064 21833 11067
rect 21600 11036 21833 11064
rect 21600 11024 21606 11036
rect 21821 11033 21833 11036
rect 21867 11033 21879 11067
rect 21821 11027 21879 11033
rect 21913 11067 21971 11073
rect 21913 11033 21925 11067
rect 21959 11064 21971 11067
rect 22002 11064 22008 11076
rect 21959 11036 22008 11064
rect 21959 11033 21971 11036
rect 21913 11027 21971 11033
rect 22002 11024 22008 11036
rect 22060 11064 22066 11076
rect 22388 11064 22416 11095
rect 22060 11036 22416 11064
rect 22060 11024 22066 11036
rect 15470 10956 15476 11008
rect 15528 10956 15534 11008
rect 1104 10906 28888 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 28888 10906
rect 1104 10832 28888 10854
rect 9214 10752 9220 10804
rect 9272 10792 9278 10804
rect 9401 10795 9459 10801
rect 9401 10792 9413 10795
rect 9272 10764 9413 10792
rect 9272 10752 9278 10764
rect 9401 10761 9413 10764
rect 9447 10761 9459 10795
rect 9401 10755 9459 10761
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 11756 10764 11836 10792
rect 11756 10752 11762 10764
rect 9766 10684 9772 10736
rect 9824 10684 9830 10736
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 11808 10733 11836 10764
rect 12894 10752 12900 10804
rect 12952 10752 12958 10804
rect 13170 10752 13176 10804
rect 13228 10752 13234 10804
rect 15746 10752 15752 10804
rect 15804 10792 15810 10804
rect 15841 10795 15899 10801
rect 15841 10792 15853 10795
rect 15804 10764 15853 10792
rect 15804 10752 15810 10764
rect 15841 10761 15853 10764
rect 15887 10761 15899 10795
rect 19518 10792 19524 10804
rect 15841 10755 15899 10761
rect 18248 10764 19524 10792
rect 11793 10727 11851 10733
rect 10192 10696 11744 10724
rect 10192 10684 10198 10696
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 9784 10656 9812 10684
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 9631 10628 11161 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 11149 10625 11161 10628
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 11330 10616 11336 10668
rect 11388 10616 11394 10668
rect 11514 10616 11520 10668
rect 11572 10616 11578 10668
rect 11716 10665 11744 10696
rect 11793 10693 11805 10727
rect 11839 10693 11851 10727
rect 11793 10687 11851 10693
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 13081 10727 13139 10733
rect 13081 10724 13093 10727
rect 12768 10696 13093 10724
rect 12768 10684 12774 10696
rect 13081 10693 13093 10696
rect 13127 10724 13139 10727
rect 14550 10724 14556 10736
rect 13127 10696 14556 10724
rect 13127 10693 13139 10696
rect 13081 10687 13139 10693
rect 14550 10684 14556 10696
rect 14608 10684 14614 10736
rect 18248 10668 18276 10764
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 19889 10795 19947 10801
rect 19889 10761 19901 10795
rect 19935 10792 19947 10795
rect 21266 10792 21272 10804
rect 19935 10764 21272 10792
rect 19935 10761 19947 10764
rect 19889 10755 19947 10761
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 24949 10795 25007 10801
rect 24949 10761 24961 10795
rect 24995 10792 25007 10795
rect 25590 10792 25596 10804
rect 24995 10764 25596 10792
rect 24995 10761 25007 10764
rect 24949 10755 25007 10761
rect 25590 10752 25596 10764
rect 25648 10752 25654 10804
rect 19610 10724 19616 10736
rect 18892 10696 19616 10724
rect 18892 10668 18920 10696
rect 19610 10684 19616 10696
rect 19668 10684 19674 10736
rect 24581 10727 24639 10733
rect 24581 10693 24593 10727
rect 24627 10724 24639 10727
rect 25130 10724 25136 10736
rect 24627 10696 25136 10724
rect 24627 10693 24639 10696
rect 24581 10687 24639 10693
rect 25130 10684 25136 10696
rect 25188 10724 25194 10736
rect 25409 10727 25467 10733
rect 25409 10724 25421 10727
rect 25188 10696 25421 10724
rect 25188 10684 25194 10696
rect 25409 10693 25421 10696
rect 25455 10693 25467 10727
rect 25409 10687 25467 10693
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11882 10616 11888 10668
rect 11940 10616 11946 10668
rect 14728 10659 14786 10665
rect 14728 10625 14740 10659
rect 14774 10656 14786 10659
rect 15194 10656 15200 10668
rect 14774 10628 15200 10656
rect 14774 10625 14786 10628
rect 14728 10619 14786 10625
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 18230 10656 18236 10668
rect 18012 10628 18236 10656
rect 18012 10616 18018 10628
rect 18230 10616 18236 10628
rect 18288 10616 18294 10668
rect 18874 10616 18880 10668
rect 18932 10616 18938 10668
rect 18984 10628 19656 10656
rect 8754 10548 8760 10600
rect 8812 10548 8818 10600
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9355 10560 9781 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 9769 10557 9781 10560
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 12069 10523 12127 10529
rect 12069 10489 12081 10523
rect 12115 10520 12127 10523
rect 12268 10520 12296 10551
rect 14458 10548 14464 10600
rect 14516 10548 14522 10600
rect 18046 10548 18052 10600
rect 18104 10548 18110 10600
rect 18138 10548 18144 10600
rect 18196 10588 18202 10600
rect 18782 10588 18788 10600
rect 18196 10560 18788 10588
rect 18196 10548 18202 10560
rect 18782 10548 18788 10560
rect 18840 10548 18846 10600
rect 18984 10588 19012 10628
rect 18892 10560 19012 10588
rect 12115 10492 12296 10520
rect 18064 10520 18092 10548
rect 18892 10520 18920 10560
rect 19426 10548 19432 10600
rect 19484 10548 19490 10600
rect 19518 10548 19524 10600
rect 19576 10548 19582 10600
rect 19628 10597 19656 10628
rect 24486 10616 24492 10668
rect 24544 10616 24550 10668
rect 24762 10616 24768 10668
rect 24820 10616 24826 10668
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 25041 10659 25099 10665
rect 25041 10656 25053 10659
rect 24912 10628 25053 10656
rect 24912 10616 24918 10628
rect 25041 10625 25053 10628
rect 25087 10625 25099 10659
rect 25041 10619 25099 10625
rect 25225 10659 25283 10665
rect 25225 10625 25237 10659
rect 25271 10656 25283 10659
rect 25958 10656 25964 10668
rect 25271 10628 25964 10656
rect 25271 10625 25283 10628
rect 25225 10619 25283 10625
rect 25958 10616 25964 10628
rect 26016 10616 26022 10668
rect 19613 10591 19671 10597
rect 19613 10557 19625 10591
rect 19659 10557 19671 10591
rect 19613 10551 19671 10557
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10557 19763 10591
rect 19705 10551 19763 10557
rect 18064 10492 18920 10520
rect 19245 10523 19303 10529
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 19245 10489 19257 10523
rect 19291 10520 19303 10523
rect 19334 10520 19340 10532
rect 19291 10492 19340 10520
rect 19291 10489 19303 10492
rect 19245 10483 19303 10489
rect 19334 10480 19340 10492
rect 19392 10520 19398 10532
rect 19720 10520 19748 10551
rect 19392 10492 19748 10520
rect 19392 10480 19398 10492
rect 10962 10412 10968 10464
rect 11020 10412 11026 10464
rect 18233 10455 18291 10461
rect 18233 10421 18245 10455
rect 18279 10452 18291 10455
rect 18414 10452 18420 10464
rect 18279 10424 18420 10452
rect 18279 10421 18291 10424
rect 18233 10415 18291 10421
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 18782 10412 18788 10464
rect 18840 10452 18846 10464
rect 19150 10452 19156 10464
rect 18840 10424 19156 10452
rect 18840 10412 18846 10424
rect 19150 10412 19156 10424
rect 19208 10452 19214 10464
rect 21358 10452 21364 10464
rect 19208 10424 21364 10452
rect 19208 10412 19214 10424
rect 21358 10412 21364 10424
rect 21416 10412 21422 10464
rect 1104 10362 28888 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 28888 10362
rect 1104 10288 28888 10310
rect 10134 10208 10140 10260
rect 10192 10208 10198 10260
rect 10597 10251 10655 10257
rect 10597 10217 10609 10251
rect 10643 10248 10655 10251
rect 11054 10248 11060 10260
rect 10643 10220 11060 10248
rect 10643 10217 10655 10220
rect 10597 10211 10655 10217
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 11333 10251 11391 10257
rect 11333 10217 11345 10251
rect 11379 10248 11391 10251
rect 11882 10248 11888 10260
rect 11379 10220 11888 10248
rect 11379 10217 11391 10220
rect 11333 10211 11391 10217
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 15194 10208 15200 10260
rect 15252 10208 15258 10260
rect 24213 10251 24271 10257
rect 24213 10217 24225 10251
rect 24259 10248 24271 10251
rect 24762 10248 24768 10260
rect 24259 10220 24768 10248
rect 24259 10217 24271 10220
rect 24213 10211 24271 10217
rect 24762 10208 24768 10220
rect 24820 10248 24826 10260
rect 24820 10220 25544 10248
rect 24820 10208 24826 10220
rect 11425 10183 11483 10189
rect 11425 10180 11437 10183
rect 11072 10152 11437 10180
rect 10778 10112 10784 10124
rect 10336 10084 10784 10112
rect 934 10004 940 10056
rect 992 10044 998 10056
rect 10336 10053 10364 10084
rect 10778 10072 10784 10084
rect 10836 10112 10842 10124
rect 11072 10121 11100 10152
rect 11425 10149 11437 10152
rect 11471 10149 11483 10183
rect 11425 10143 11483 10149
rect 17512 10152 19012 10180
rect 11057 10115 11115 10121
rect 11057 10112 11069 10115
rect 10836 10084 11069 10112
rect 10836 10072 10842 10084
rect 11057 10081 11069 10084
rect 11103 10081 11115 10115
rect 11057 10075 11115 10081
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 11514 10112 11520 10124
rect 11195 10084 11520 10112
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 17512 10121 17540 10152
rect 17497 10115 17555 10121
rect 17497 10081 17509 10115
rect 17543 10081 17555 10115
rect 17497 10075 17555 10081
rect 18414 10072 18420 10124
rect 18472 10072 18478 10124
rect 18506 10072 18512 10124
rect 18564 10072 18570 10124
rect 18877 10115 18935 10121
rect 18877 10112 18889 10115
rect 18616 10084 18889 10112
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 992 10016 1409 10044
rect 992 10004 998 10016
rect 1397 10013 1409 10016
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12124 10016 12817 10044
rect 12124 10004 12130 10016
rect 12805 10013 12817 10016
rect 12851 10044 12863 10047
rect 14458 10044 14464 10056
rect 12851 10016 14464 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 15010 10004 15016 10056
rect 15068 10004 15074 10056
rect 15197 10047 15255 10053
rect 15197 10013 15209 10047
rect 15243 10044 15255 10047
rect 15470 10044 15476 10056
rect 15243 10016 15476 10044
rect 15243 10013 15255 10016
rect 15197 10007 15255 10013
rect 15470 10004 15476 10016
rect 15528 10004 15534 10056
rect 17681 10047 17739 10053
rect 17681 10013 17693 10047
rect 17727 10044 17739 10047
rect 18138 10044 18144 10056
rect 17727 10016 18144 10044
rect 17727 10013 17739 10016
rect 17681 10007 17739 10013
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18616 10044 18644 10084
rect 18877 10081 18889 10084
rect 18923 10081 18935 10115
rect 18877 10075 18935 10081
rect 18380 10016 18644 10044
rect 18785 10047 18843 10053
rect 18380 10004 18386 10016
rect 18785 10013 18797 10047
rect 18831 10044 18843 10047
rect 18984 10044 19012 10152
rect 21358 10140 21364 10192
rect 21416 10180 21422 10192
rect 24854 10180 24860 10192
rect 21416 10152 24860 10180
rect 21416 10140 21422 10152
rect 19334 10072 19340 10124
rect 19392 10072 19398 10124
rect 19058 10044 19064 10056
rect 18831 10016 19064 10044
rect 18831 10013 18843 10016
rect 18785 10007 18843 10013
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 24044 10053 24072 10152
rect 24854 10140 24860 10152
rect 24912 10140 24918 10192
rect 25130 10140 25136 10192
rect 25188 10140 25194 10192
rect 24486 10072 24492 10124
rect 24544 10072 24550 10124
rect 25516 10121 25544 10220
rect 25590 10208 25596 10260
rect 25648 10248 25654 10260
rect 25685 10251 25743 10257
rect 25685 10248 25697 10251
rect 25648 10220 25697 10248
rect 25648 10208 25654 10220
rect 25685 10217 25697 10220
rect 25731 10248 25743 10251
rect 26786 10248 26792 10260
rect 25731 10220 26792 10248
rect 25731 10217 25743 10220
rect 25685 10211 25743 10217
rect 26786 10208 26792 10220
rect 26844 10208 26850 10260
rect 25041 10115 25099 10121
rect 25041 10081 25053 10115
rect 25087 10081 25099 10115
rect 25041 10075 25099 10081
rect 25501 10115 25559 10121
rect 25501 10081 25513 10115
rect 25547 10081 25559 10115
rect 25501 10075 25559 10081
rect 25608 10084 26004 10112
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 23937 10047 23995 10053
rect 23937 10013 23949 10047
rect 23983 10013 23995 10047
rect 23937 10007 23995 10013
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10013 24087 10047
rect 24029 10007 24087 10013
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10044 24639 10047
rect 25056 10044 25084 10075
rect 24627 10016 25084 10044
rect 24627 10013 24639 10016
rect 24581 10007 24639 10013
rect 10594 9936 10600 9988
rect 10652 9936 10658 9988
rect 10781 9979 10839 9985
rect 10781 9945 10793 9979
rect 10827 9976 10839 9979
rect 10962 9976 10968 9988
rect 10827 9948 10968 9976
rect 10827 9945 10839 9948
rect 10781 9939 10839 9945
rect 10962 9936 10968 9948
rect 11020 9976 11026 9988
rect 12538 9979 12596 9985
rect 12538 9976 12550 9979
rect 11020 9948 12550 9976
rect 11020 9936 11026 9948
rect 12538 9945 12550 9948
rect 12584 9945 12596 9979
rect 12538 9939 12596 9945
rect 17865 9979 17923 9985
rect 17865 9945 17877 9979
rect 17911 9976 17923 9979
rect 18598 9976 18604 9988
rect 17911 9948 18604 9976
rect 17911 9945 17923 9948
rect 17865 9939 17923 9945
rect 18598 9936 18604 9948
rect 18656 9936 18662 9988
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 19444 9976 19472 10007
rect 19392 9948 19472 9976
rect 23952 9976 23980 10007
rect 25608 9976 25636 10084
rect 25976 10056 26004 10084
rect 25869 10047 25927 10053
rect 25869 10013 25881 10047
rect 25915 10013 25927 10047
rect 25869 10007 25927 10013
rect 23952 9948 25636 9976
rect 25884 9976 25912 10007
rect 25958 10004 25964 10056
rect 26016 10004 26022 10056
rect 28350 9976 28356 9988
rect 25884 9948 28356 9976
rect 19392 9936 19398 9948
rect 28350 9936 28356 9948
rect 28408 9936 28414 9988
rect 10873 9911 10931 9917
rect 10873 9877 10885 9911
rect 10919 9908 10931 9911
rect 11054 9908 11060 9920
rect 10919 9880 11060 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 11054 9868 11060 9880
rect 11112 9908 11118 9920
rect 11514 9908 11520 9920
rect 11112 9880 11520 9908
rect 11112 9868 11118 9880
rect 11514 9868 11520 9880
rect 11572 9868 11578 9920
rect 17954 9868 17960 9920
rect 18012 9868 18018 9920
rect 18138 9868 18144 9920
rect 18196 9908 18202 9920
rect 18506 9908 18512 9920
rect 18196 9880 18512 9908
rect 18196 9868 18202 9880
rect 18506 9868 18512 9880
rect 18564 9908 18570 9920
rect 19518 9908 19524 9920
rect 18564 9880 19524 9908
rect 18564 9868 18570 9880
rect 19518 9868 19524 9880
rect 19576 9868 19582 9920
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 19797 9911 19855 9917
rect 19797 9908 19809 9911
rect 19760 9880 19809 9908
rect 19760 9868 19766 9880
rect 19797 9877 19809 9880
rect 19843 9877 19855 9911
rect 19797 9871 19855 9877
rect 24946 9868 24952 9920
rect 25004 9868 25010 9920
rect 25222 9868 25228 9920
rect 25280 9908 25286 9920
rect 26053 9911 26111 9917
rect 26053 9908 26065 9911
rect 25280 9880 26065 9908
rect 25280 9868 25286 9880
rect 26053 9877 26065 9880
rect 26099 9877 26111 9911
rect 26053 9871 26111 9877
rect 1104 9818 28888 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 28888 9818
rect 1104 9744 28888 9766
rect 10321 9707 10379 9713
rect 10321 9673 10333 9707
rect 10367 9704 10379 9707
rect 10410 9704 10416 9716
rect 10367 9676 10416 9704
rect 10367 9673 10379 9676
rect 10321 9667 10379 9673
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 10505 9707 10563 9713
rect 10505 9673 10517 9707
rect 10551 9704 10563 9707
rect 10686 9704 10692 9716
rect 10551 9676 10692 9704
rect 10551 9673 10563 9676
rect 10505 9667 10563 9673
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11514 9664 11520 9716
rect 11572 9664 11578 9716
rect 16022 9704 16028 9716
rect 15304 9676 16028 9704
rect 9306 9636 9312 9648
rect 7208 9608 9312 9636
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 7208 9577 7236 9608
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 9950 9596 9956 9648
rect 10008 9636 10014 9648
rect 10229 9639 10287 9645
rect 10229 9636 10241 9639
rect 10008 9608 10241 9636
rect 10008 9596 10014 9608
rect 10229 9605 10241 9608
rect 10275 9605 10287 9639
rect 10229 9599 10287 9605
rect 14550 9596 14556 9648
rect 14608 9596 14614 9648
rect 15010 9596 15016 9648
rect 15068 9596 15074 9648
rect 15194 9596 15200 9648
rect 15252 9596 15258 9648
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 5868 9540 7205 9568
rect 5868 9528 5874 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 7449 9571 7507 9577
rect 7449 9568 7461 9571
rect 7340 9540 7461 9568
rect 7340 9528 7346 9540
rect 7449 9537 7461 9540
rect 7495 9537 7507 9571
rect 7449 9531 7507 9537
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 9766 9568 9772 9580
rect 9723 9540 9772 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 10778 9528 10784 9580
rect 10836 9528 10842 9580
rect 12158 9528 12164 9580
rect 12216 9568 12222 9580
rect 12630 9571 12688 9577
rect 12630 9568 12642 9571
rect 12216 9540 12642 9568
rect 12216 9528 12222 9540
rect 12630 9537 12642 9540
rect 12676 9537 12688 9571
rect 12630 9531 12688 9537
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9568 14703 9571
rect 15028 9568 15056 9596
rect 15304 9577 15332 9676
rect 16022 9664 16028 9676
rect 16080 9704 16086 9716
rect 18138 9704 18144 9716
rect 16080 9676 18144 9704
rect 16080 9664 16086 9676
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 18230 9664 18236 9716
rect 18288 9704 18294 9716
rect 18417 9707 18475 9713
rect 18417 9704 18429 9707
rect 18288 9676 18429 9704
rect 18288 9664 18294 9676
rect 18417 9673 18429 9676
rect 18463 9673 18475 9707
rect 18417 9667 18475 9673
rect 19426 9664 19432 9716
rect 19484 9664 19490 9716
rect 24946 9664 24952 9716
rect 25004 9704 25010 9716
rect 25041 9707 25099 9713
rect 25041 9704 25053 9707
rect 25004 9676 25053 9704
rect 25004 9664 25010 9676
rect 25041 9673 25053 9676
rect 25087 9673 25099 9707
rect 25041 9667 25099 9673
rect 18785 9639 18843 9645
rect 18785 9605 18797 9639
rect 18831 9636 18843 9639
rect 19334 9636 19340 9648
rect 18831 9608 19340 9636
rect 18831 9605 18843 9608
rect 18785 9599 18843 9605
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 24029 9639 24087 9645
rect 24029 9636 24041 9639
rect 23768 9608 24041 9636
rect 14691 9540 15056 9568
rect 15289 9571 15347 9577
rect 14691 9537 14703 9540
rect 14645 9531 14703 9537
rect 15289 9537 15301 9571
rect 15335 9568 15347 9571
rect 15378 9568 15384 9580
rect 15335 9540 15384 9568
rect 15335 9537 15347 9540
rect 15289 9531 15347 9537
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 18046 9528 18052 9580
rect 18104 9568 18110 9580
rect 18325 9571 18383 9577
rect 18325 9568 18337 9571
rect 18104 9540 18337 9568
rect 18104 9528 18110 9540
rect 18325 9537 18337 9540
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 18598 9528 18604 9580
rect 18656 9528 18662 9580
rect 19058 9528 19064 9580
rect 19116 9528 19122 9580
rect 19150 9528 19156 9580
rect 19208 9568 19214 9580
rect 19245 9571 19303 9577
rect 19245 9568 19257 9571
rect 19208 9540 19257 9568
rect 19208 9528 19214 9540
rect 19245 9537 19257 9540
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 21542 9568 21548 9580
rect 21315 9540 21548 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 21542 9528 21548 9540
rect 21600 9528 21606 9580
rect 22002 9568 22008 9580
rect 21652 9540 22008 9568
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 9456 9472 9505 9500
rect 9456 9460 9462 9472
rect 9493 9469 9505 9472
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 14458 9500 14464 9512
rect 12943 9472 14464 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9500 19027 9503
rect 20070 9500 20076 9512
rect 19015 9472 20076 9500
rect 19015 9469 19027 9472
rect 18969 9463 19027 9469
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 21174 9460 21180 9512
rect 21232 9460 21238 9512
rect 21652 9509 21680 9540
rect 22002 9528 22008 9540
rect 22060 9528 22066 9580
rect 23768 9577 23796 9608
rect 24029 9605 24041 9608
rect 24075 9605 24087 9639
rect 24029 9599 24087 9605
rect 24397 9639 24455 9645
rect 24397 9605 24409 9639
rect 24443 9636 24455 9639
rect 25406 9636 25412 9648
rect 24443 9608 25412 9636
rect 24443 9605 24455 9608
rect 24397 9599 24455 9605
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 25590 9596 25596 9648
rect 25648 9596 25654 9648
rect 23753 9571 23811 9577
rect 23753 9537 23765 9571
rect 23799 9537 23811 9571
rect 23753 9531 23811 9537
rect 23937 9571 23995 9577
rect 23937 9537 23949 9571
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 21637 9503 21695 9509
rect 21637 9469 21649 9503
rect 21683 9469 21695 9503
rect 21637 9463 21695 9469
rect 21910 9460 21916 9512
rect 21968 9460 21974 9512
rect 23768 9500 23796 9531
rect 22066 9472 23796 9500
rect 23952 9500 23980 9531
rect 24578 9528 24584 9580
rect 24636 9568 24642 9580
rect 24949 9571 25007 9577
rect 24636 9540 24716 9568
rect 24636 9528 24642 9540
rect 24688 9500 24716 9540
rect 24949 9537 24961 9571
rect 24995 9568 25007 9571
rect 25222 9568 25228 9580
rect 24995 9540 25228 9568
rect 24995 9537 25007 9540
rect 24949 9531 25007 9537
rect 25222 9528 25228 9540
rect 25280 9528 25286 9580
rect 25133 9503 25191 9509
rect 25133 9500 25145 9503
rect 23952 9472 24624 9500
rect 24688 9472 25145 9500
rect 22066 9444 22094 9472
rect 8573 9435 8631 9441
rect 8573 9401 8585 9435
rect 8619 9432 8631 9435
rect 8754 9432 8760 9444
rect 8619 9404 8760 9432
rect 8619 9401 8631 9404
rect 8573 9395 8631 9401
rect 8754 9392 8760 9404
rect 8812 9432 8818 9444
rect 9953 9435 10011 9441
rect 9953 9432 9965 9435
rect 8812 9404 9965 9432
rect 8812 9392 8818 9404
rect 9953 9401 9965 9404
rect 9999 9432 10011 9435
rect 10778 9432 10784 9444
rect 9999 9404 10784 9432
rect 9999 9401 10011 9404
rect 9953 9395 10011 9401
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 20714 9392 20720 9444
rect 20772 9432 20778 9444
rect 22002 9432 22008 9444
rect 20772 9404 22008 9432
rect 20772 9392 20778 9404
rect 22002 9392 22008 9404
rect 22060 9404 22094 9444
rect 24596 9441 24624 9472
rect 25133 9469 25145 9472
rect 25179 9469 25191 9503
rect 25133 9463 25191 9469
rect 24581 9435 24639 9441
rect 22060 9392 22066 9404
rect 24581 9401 24593 9435
rect 24627 9401 24639 9435
rect 24581 9395 24639 9401
rect 9858 9324 9864 9376
rect 9916 9324 9922 9376
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 11204 9336 11345 9364
rect 11204 9324 11210 9336
rect 11333 9333 11345 9336
rect 11379 9333 11391 9367
rect 11333 9327 11391 9333
rect 14918 9324 14924 9376
rect 14976 9364 14982 9376
rect 15013 9367 15071 9373
rect 15013 9364 15025 9367
rect 14976 9336 15025 9364
rect 14976 9324 14982 9336
rect 15013 9333 15025 9336
rect 15059 9333 15071 9367
rect 15013 9327 15071 9333
rect 22281 9367 22339 9373
rect 22281 9333 22293 9367
rect 22327 9364 22339 9367
rect 22462 9364 22468 9376
rect 22327 9336 22468 9364
rect 22327 9333 22339 9336
rect 22281 9327 22339 9333
rect 22462 9324 22468 9336
rect 22520 9324 22526 9376
rect 23934 9324 23940 9376
rect 23992 9324 23998 9376
rect 1104 9274 28888 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 28888 9274
rect 1104 9200 28888 9222
rect 9398 9120 9404 9172
rect 9456 9120 9462 9172
rect 10505 9163 10563 9169
rect 10505 9129 10517 9163
rect 10551 9129 10563 9163
rect 10505 9123 10563 9129
rect 7193 9095 7251 9101
rect 7193 9061 7205 9095
rect 7239 9092 7251 9095
rect 10134 9092 10140 9104
rect 7239 9064 10140 9092
rect 7239 9061 7251 9064
rect 7193 9055 7251 9061
rect 5810 8984 5816 9036
rect 5868 8984 5874 9036
rect 8036 9033 8064 9064
rect 10134 9052 10140 9064
rect 10192 9092 10198 9104
rect 10520 9092 10548 9123
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 10965 9163 11023 9169
rect 10965 9160 10977 9163
rect 10652 9132 10977 9160
rect 10652 9120 10658 9132
rect 10965 9129 10977 9132
rect 11011 9129 11023 9163
rect 10965 9123 11023 9129
rect 12158 9120 12164 9172
rect 12216 9120 12222 9172
rect 15286 9120 15292 9172
rect 15344 9160 15350 9172
rect 15565 9163 15623 9169
rect 15565 9160 15577 9163
rect 15344 9132 15577 9160
rect 15344 9120 15350 9132
rect 15565 9129 15577 9132
rect 15611 9129 15623 9163
rect 15565 9123 15623 9129
rect 21729 9163 21787 9169
rect 21729 9129 21741 9163
rect 21775 9160 21787 9163
rect 22370 9160 22376 9172
rect 21775 9132 22376 9160
rect 21775 9129 21787 9132
rect 21729 9123 21787 9129
rect 10192 9064 10548 9092
rect 10192 9052 10198 9064
rect 19518 9052 19524 9104
rect 19576 9092 19582 9104
rect 21744 9092 21772 9123
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 25777 9163 25835 9169
rect 25777 9129 25789 9163
rect 25823 9160 25835 9163
rect 25958 9160 25964 9172
rect 25823 9132 25964 9160
rect 25823 9129 25835 9132
rect 25777 9123 25835 9129
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 19576 9064 21772 9092
rect 19576 9052 19582 9064
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 10594 8984 10600 9036
rect 10652 8984 10658 9036
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 11020 8996 12541 9024
rect 11020 8984 11026 8996
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 10008 8928 10517 8956
rect 10008 8916 10014 8928
rect 10505 8925 10517 8928
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 10778 8916 10784 8968
rect 10836 8916 10842 8968
rect 11992 8965 12020 8996
rect 12529 8993 12541 8996
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 19702 8984 19708 9036
rect 19760 8984 19766 9036
rect 19904 9033 19932 9064
rect 21910 9052 21916 9104
rect 21968 9092 21974 9104
rect 22189 9095 22247 9101
rect 22189 9092 22201 9095
rect 21968 9064 22201 9092
rect 21968 9052 21974 9064
rect 22189 9061 22201 9064
rect 22235 9061 22247 9095
rect 22189 9055 22247 9061
rect 19889 9027 19947 9033
rect 19889 8993 19901 9027
rect 19935 8993 19947 9027
rect 19889 8987 19947 8993
rect 21542 8984 21548 9036
rect 21600 9024 21606 9036
rect 21637 9027 21695 9033
rect 21637 9024 21649 9027
rect 21600 8996 21649 9024
rect 21600 8984 21606 8996
rect 21637 8993 21649 8996
rect 21683 8993 21695 9027
rect 21637 8987 21695 8993
rect 21818 8984 21824 9036
rect 21876 9024 21882 9036
rect 24397 9027 24455 9033
rect 24397 9024 24409 9027
rect 21876 8996 24409 9024
rect 21876 8984 21882 8996
rect 24397 8993 24409 8996
rect 24443 8993 24455 9027
rect 24397 8987 24455 8993
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8956 11759 8959
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11747 8928 11805 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 11793 8925 11805 8928
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8925 12035 8959
rect 11977 8919 12035 8925
rect 14185 8959 14243 8965
rect 14185 8925 14197 8959
rect 14231 8956 14243 8959
rect 14274 8956 14280 8968
rect 14231 8928 14280 8956
rect 14231 8925 14243 8928
rect 14185 8919 14243 8925
rect 5626 8848 5632 8900
rect 5684 8888 5690 8900
rect 6058 8891 6116 8897
rect 6058 8888 6070 8891
rect 5684 8860 6070 8888
rect 5684 8848 5690 8860
rect 6058 8857 6070 8860
rect 6104 8857 6116 8891
rect 6058 8851 6116 8857
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 11072 8888 11100 8919
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 15010 8916 15016 8968
rect 15068 8956 15074 8968
rect 17221 8959 17279 8965
rect 17221 8956 17233 8959
rect 15068 8928 17233 8956
rect 15068 8916 15074 8928
rect 17221 8925 17233 8928
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 17405 8959 17463 8965
rect 17405 8925 17417 8959
rect 17451 8956 17463 8959
rect 17954 8956 17960 8968
rect 17451 8928 17960 8956
rect 17451 8925 17463 8928
rect 17405 8919 17463 8925
rect 10468 8860 11100 8888
rect 10468 8848 10474 8860
rect 12342 8848 12348 8900
rect 12400 8848 12406 8900
rect 14452 8891 14510 8897
rect 14452 8857 14464 8891
rect 14498 8888 14510 8891
rect 14734 8888 14740 8900
rect 14498 8860 14740 8888
rect 14498 8857 14510 8860
rect 14452 8851 14510 8857
rect 14734 8848 14740 8860
rect 14792 8848 14798 8900
rect 17236 8888 17264 8919
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 19610 8916 19616 8968
rect 19668 8916 19674 8968
rect 20070 8916 20076 8968
rect 20128 8916 20134 8968
rect 21910 8916 21916 8968
rect 21968 8916 21974 8968
rect 22462 8916 22468 8968
rect 22520 8916 22526 8968
rect 23934 8916 23940 8968
rect 23992 8956 23998 8968
rect 24653 8959 24711 8965
rect 24653 8956 24665 8959
rect 23992 8928 24665 8956
rect 23992 8916 23998 8928
rect 24653 8925 24665 8928
rect 24699 8925 24711 8959
rect 24653 8919 24711 8925
rect 18690 8888 18696 8900
rect 17236 8860 18696 8888
rect 18690 8848 18696 8860
rect 18748 8848 18754 8900
rect 19628 8888 19656 8916
rect 20165 8891 20223 8897
rect 20165 8888 20177 8891
rect 19628 8860 20177 8888
rect 20165 8857 20177 8860
rect 20211 8857 20223 8891
rect 20165 8851 20223 8857
rect 22002 8848 22008 8900
rect 22060 8888 22066 8900
rect 22189 8891 22247 8897
rect 22189 8888 22201 8891
rect 22060 8860 22201 8888
rect 22060 8848 22066 8860
rect 22189 8857 22201 8860
rect 22235 8857 22247 8891
rect 22189 8851 22247 8857
rect 7469 8823 7527 8829
rect 7469 8789 7481 8823
rect 7515 8820 7527 8823
rect 7558 8820 7564 8832
rect 7515 8792 7564 8820
rect 7515 8789 7527 8792
rect 7469 8783 7527 8789
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 17313 8823 17371 8829
rect 17313 8820 17325 8823
rect 17276 8792 17325 8820
rect 17276 8780 17282 8792
rect 17313 8789 17325 8792
rect 17359 8789 17371 8823
rect 17313 8783 17371 8789
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 19245 8823 19303 8829
rect 19245 8820 19257 8823
rect 18932 8792 19257 8820
rect 18932 8780 18938 8792
rect 19245 8789 19257 8792
rect 19291 8789 19303 8823
rect 19245 8783 19303 8789
rect 22094 8780 22100 8832
rect 22152 8780 22158 8832
rect 22370 8780 22376 8832
rect 22428 8820 22434 8832
rect 24578 8820 24584 8832
rect 22428 8792 24584 8820
rect 22428 8780 22434 8792
rect 24578 8780 24584 8792
rect 24636 8780 24642 8832
rect 1104 8730 28888 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 28888 8730
rect 1104 8656 28888 8678
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 7282 8576 7288 8628
rect 7340 8576 7346 8628
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 9824 8588 10364 8616
rect 9824 8576 9830 8588
rect 7834 8548 7840 8560
rect 5368 8520 7840 8548
rect 5368 8489 5396 8520
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5442 8440 5448 8492
rect 5500 8440 5506 8492
rect 7484 8489 7512 8520
rect 7834 8508 7840 8520
rect 7892 8508 7898 8560
rect 9576 8551 9634 8557
rect 9576 8517 9588 8551
rect 9622 8548 9634 8551
rect 9858 8548 9864 8560
rect 9622 8520 9864 8548
rect 9622 8517 9634 8520
rect 9576 8511 9634 8517
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 10336 8548 10364 8588
rect 10410 8576 10416 8628
rect 10468 8616 10474 8628
rect 10689 8619 10747 8625
rect 10689 8616 10701 8619
rect 10468 8588 10701 8616
rect 10468 8576 10474 8588
rect 10689 8585 10701 8588
rect 10735 8585 10747 8619
rect 10689 8579 10747 8585
rect 14734 8576 14740 8628
rect 14792 8576 14798 8628
rect 18325 8619 18383 8625
rect 18325 8585 18337 8619
rect 18371 8616 18383 8619
rect 19058 8616 19064 8628
rect 18371 8588 19064 8616
rect 18371 8585 18383 8588
rect 18325 8579 18383 8585
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 21542 8576 21548 8628
rect 21600 8616 21606 8628
rect 23201 8619 23259 8625
rect 23201 8616 23213 8619
rect 21600 8588 23213 8616
rect 21600 8576 21606 8588
rect 23201 8585 23213 8588
rect 23247 8585 23259 8619
rect 23201 8579 23259 8585
rect 28350 8576 28356 8628
rect 28408 8576 28414 8628
rect 11885 8551 11943 8557
rect 10336 8520 10916 8548
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 7558 8440 7564 8492
rect 7616 8440 7622 8492
rect 7852 8480 7880 8508
rect 10888 8480 10916 8520
rect 11885 8517 11897 8551
rect 11931 8548 11943 8551
rect 13170 8548 13176 8560
rect 11931 8520 13176 8548
rect 11931 8517 11943 8520
rect 11885 8511 11943 8517
rect 13170 8508 13176 8520
rect 13228 8508 13234 8560
rect 14458 8508 14464 8560
rect 14516 8548 14522 8560
rect 22094 8557 22100 8560
rect 14516 8520 19288 8548
rect 14516 8508 14522 8520
rect 10962 8480 10968 8492
rect 7852 8452 10364 8480
rect 10888 8452 10968 8480
rect 9306 8372 9312 8424
rect 9364 8372 9370 8424
rect 10336 8412 10364 8452
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 11146 8440 11152 8492
rect 11204 8440 11210 8492
rect 14918 8440 14924 8492
rect 14976 8440 14982 8492
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 15286 8480 15292 8492
rect 15243 8452 15292 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 16960 8489 16988 8520
rect 19260 8492 19288 8520
rect 22088 8511 22100 8557
rect 22152 8548 22158 8560
rect 22152 8520 22188 8548
rect 22094 8508 22100 8511
rect 22152 8508 22158 8520
rect 17218 8489 17224 8492
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 17212 8480 17224 8489
rect 17179 8452 17224 8480
rect 16945 8443 17003 8449
rect 17212 8443 17224 8452
rect 17218 8440 17224 8443
rect 17276 8440 17282 8492
rect 18690 8440 18696 8492
rect 18748 8440 18754 8492
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 19242 8440 19248 8492
rect 19300 8480 19306 8492
rect 21818 8480 21824 8492
rect 19300 8452 21824 8480
rect 19300 8440 19306 8452
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 28534 8440 28540 8492
rect 28592 8440 28598 8492
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 10336 8384 11713 8412
rect 11701 8381 11713 8384
rect 11747 8412 11759 8415
rect 12342 8412 12348 8424
rect 11747 8384 12348 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 15105 8415 15163 8421
rect 15105 8381 15117 8415
rect 15151 8412 15163 8415
rect 15378 8412 15384 8424
rect 15151 8384 15384 8412
rect 15151 8381 15163 8384
rect 15105 8375 15163 8381
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 18708 8412 18736 8440
rect 20714 8412 20720 8424
rect 18708 8384 20720 8412
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 18877 8347 18935 8353
rect 18877 8313 18889 8347
rect 18923 8344 18935 8347
rect 19334 8344 19340 8356
rect 18923 8316 19340 8344
rect 18923 8313 18935 8316
rect 18877 8307 18935 8313
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 10778 8236 10784 8288
rect 10836 8236 10842 8288
rect 1104 8186 28888 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 28888 8186
rect 1104 8112 28888 8134
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9950 8072 9956 8084
rect 8987 8044 9956 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 20625 8075 20683 8081
rect 20625 8072 20637 8075
rect 20220 8044 20637 8072
rect 20220 8032 20226 8044
rect 20625 8041 20637 8044
rect 20671 8041 20683 8075
rect 20625 8035 20683 8041
rect 19242 7896 19248 7948
rect 19300 7896 19306 7948
rect 9306 7828 9312 7880
rect 9364 7868 9370 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 9364 7840 10333 7868
rect 9364 7828 9370 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19501 7871 19559 7877
rect 19501 7868 19513 7871
rect 19392 7840 19513 7868
rect 19392 7828 19398 7840
rect 19501 7837 19513 7840
rect 19547 7837 19559 7871
rect 19501 7831 19559 7837
rect 10076 7803 10134 7809
rect 10076 7769 10088 7803
rect 10122 7800 10134 7803
rect 10778 7800 10784 7812
rect 10122 7772 10784 7800
rect 10122 7769 10134 7772
rect 10076 7763 10134 7769
rect 10778 7760 10784 7772
rect 10836 7760 10842 7812
rect 1104 7642 28888 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 28888 7642
rect 1104 7568 28888 7590
rect 1104 7098 28888 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 28888 7098
rect 1104 7024 28888 7046
rect 1104 6554 28888 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 28888 6554
rect 1104 6480 28888 6502
rect 1104 6010 28888 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 28888 6010
rect 1104 5936 28888 5958
rect 1104 5466 28888 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 28888 5466
rect 1104 5392 28888 5414
rect 1104 4922 28888 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 28888 4922
rect 1104 4848 28888 4870
rect 1104 4378 28888 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 28888 3290
rect 1104 3216 28888 3238
rect 1104 2746 28888 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 28888 2746
rect 1104 2672 28888 2694
rect 5442 2592 5448 2644
rect 5500 2592 5506 2644
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 1104 2202 28888 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 7104 47132 7156 47184
rect 6552 47039 6604 47048
rect 6552 47005 6561 47039
rect 6561 47005 6595 47039
rect 6595 47005 6604 47039
rect 6552 46996 6604 47005
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 7104 45475 7156 45484
rect 7104 45441 7113 45475
rect 7113 45441 7147 45475
rect 7147 45441 7156 45475
rect 7104 45432 7156 45441
rect 8208 45364 8260 45416
rect 12348 45432 12400 45484
rect 12072 45407 12124 45416
rect 12072 45373 12081 45407
rect 12081 45373 12115 45407
rect 12115 45373 12124 45407
rect 12072 45364 12124 45373
rect 12256 45296 12308 45348
rect 7288 45271 7340 45280
rect 7288 45237 7297 45271
rect 7297 45237 7331 45271
rect 7331 45237 7340 45271
rect 7288 45228 7340 45237
rect 12164 45271 12216 45280
rect 12164 45237 12173 45271
rect 12173 45237 12207 45271
rect 12207 45237 12216 45271
rect 12164 45228 12216 45237
rect 12440 45271 12492 45280
rect 12440 45237 12449 45271
rect 12449 45237 12483 45271
rect 12483 45237 12492 45271
rect 12440 45228 12492 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 12072 45024 12124 45076
rect 9588 44888 9640 44940
rect 12532 44931 12584 44940
rect 12532 44897 12541 44931
rect 12541 44897 12575 44931
rect 12575 44897 12584 44931
rect 12532 44888 12584 44897
rect 13544 44888 13596 44940
rect 7288 44752 7340 44804
rect 12256 44863 12308 44872
rect 12256 44829 12265 44863
rect 12265 44829 12299 44863
rect 12299 44829 12308 44863
rect 12256 44820 12308 44829
rect 13820 44820 13872 44872
rect 8944 44727 8996 44736
rect 8944 44693 8953 44727
rect 8953 44693 8987 44727
rect 8987 44693 8996 44727
rect 8944 44684 8996 44693
rect 11520 44752 11572 44804
rect 12164 44752 12216 44804
rect 12624 44752 12676 44804
rect 14464 44752 14516 44804
rect 11888 44684 11940 44736
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 12256 44480 12308 44532
rect 13268 44480 13320 44532
rect 8944 44412 8996 44464
rect 12532 44412 12584 44464
rect 9588 44344 9640 44396
rect 9772 44319 9824 44328
rect 9772 44285 9781 44319
rect 9781 44285 9815 44319
rect 9815 44285 9824 44319
rect 9772 44276 9824 44285
rect 11704 44344 11756 44396
rect 12072 44344 12124 44396
rect 13176 44344 13228 44396
rect 13544 44344 13596 44396
rect 14464 44344 14516 44396
rect 8576 44183 8628 44192
rect 8576 44149 8585 44183
rect 8585 44149 8619 44183
rect 8619 44149 8628 44183
rect 8576 44140 8628 44149
rect 11796 44183 11848 44192
rect 11796 44149 11805 44183
rect 11805 44149 11839 44183
rect 11839 44149 11848 44183
rect 11796 44140 11848 44149
rect 12716 44140 12768 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 9588 43936 9640 43988
rect 9864 43936 9916 43988
rect 11520 43979 11572 43988
rect 11520 43945 11529 43979
rect 11529 43945 11563 43979
rect 11563 43945 11572 43979
rect 11520 43936 11572 43945
rect 12440 43936 12492 43988
rect 13176 43979 13228 43988
rect 13176 43945 13185 43979
rect 13185 43945 13219 43979
rect 13219 43945 13228 43979
rect 13176 43936 13228 43945
rect 13268 43979 13320 43988
rect 13268 43945 13277 43979
rect 13277 43945 13311 43979
rect 13311 43945 13320 43979
rect 13268 43936 13320 43945
rect 11888 43843 11940 43852
rect 11888 43809 11897 43843
rect 11897 43809 11931 43843
rect 11931 43809 11940 43843
rect 11888 43800 11940 43809
rect 12348 43800 12400 43852
rect 8576 43732 8628 43784
rect 11704 43775 11756 43784
rect 11704 43741 11713 43775
rect 11713 43741 11747 43775
rect 11747 43741 11756 43775
rect 11704 43732 11756 43741
rect 12992 43868 13044 43920
rect 12716 43800 12768 43852
rect 12624 43775 12676 43784
rect 12624 43741 12633 43775
rect 12633 43741 12667 43775
rect 12667 43741 12676 43775
rect 12624 43732 12676 43741
rect 12992 43775 13044 43784
rect 12992 43741 13001 43775
rect 13001 43741 13035 43775
rect 13035 43741 13044 43775
rect 12992 43732 13044 43741
rect 13176 43732 13228 43784
rect 13820 43732 13872 43784
rect 14648 43775 14700 43784
rect 14648 43741 14657 43775
rect 14657 43741 14691 43775
rect 14691 43741 14700 43775
rect 14648 43732 14700 43741
rect 12164 43596 12216 43648
rect 12624 43596 12676 43648
rect 12808 43596 12860 43648
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 11704 43392 11756 43444
rect 13360 43392 13412 43444
rect 13820 43392 13872 43444
rect 14648 43392 14700 43444
rect 11704 43299 11756 43308
rect 11704 43265 11710 43299
rect 11710 43265 11744 43299
rect 11744 43265 11756 43299
rect 11704 43256 11756 43265
rect 11796 43299 11848 43308
rect 11796 43265 11805 43299
rect 11805 43265 11839 43299
rect 11839 43265 11848 43299
rect 11796 43256 11848 43265
rect 12532 43256 12584 43308
rect 12992 43299 13044 43308
rect 12992 43265 13026 43299
rect 13026 43265 13044 43299
rect 12992 43256 13044 43265
rect 22836 43324 22888 43376
rect 20168 43299 20220 43308
rect 20168 43265 20202 43299
rect 20202 43265 20220 43299
rect 20168 43256 20220 43265
rect 12440 43188 12492 43240
rect 11336 43052 11388 43104
rect 12716 43052 12768 43104
rect 21272 43095 21324 43104
rect 21272 43061 21281 43095
rect 21281 43061 21315 43095
rect 21315 43061 21324 43095
rect 21272 43052 21324 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 12440 42891 12492 42900
rect 12440 42857 12449 42891
rect 12449 42857 12483 42891
rect 12483 42857 12492 42891
rect 12440 42848 12492 42857
rect 12992 42848 13044 42900
rect 9588 42712 9640 42764
rect 21272 42712 21324 42764
rect 11336 42687 11388 42696
rect 11336 42653 11370 42687
rect 11370 42653 11388 42687
rect 11336 42644 11388 42653
rect 12624 42644 12676 42696
rect 12808 42687 12860 42696
rect 12808 42653 12817 42687
rect 12817 42653 12851 42687
rect 12851 42653 12860 42687
rect 12808 42644 12860 42653
rect 13268 42687 13320 42696
rect 13268 42653 13277 42687
rect 13277 42653 13311 42687
rect 13311 42653 13320 42687
rect 13268 42644 13320 42653
rect 12716 42508 12768 42560
rect 12992 42551 13044 42560
rect 12992 42517 13001 42551
rect 13001 42517 13035 42551
rect 13035 42517 13044 42551
rect 12992 42508 13044 42517
rect 20812 42508 20864 42560
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 12992 42168 13044 42220
rect 12624 41964 12676 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 20168 41803 20220 41812
rect 20168 41769 20177 41803
rect 20177 41769 20211 41803
rect 20211 41769 20220 41803
rect 20168 41760 20220 41769
rect 17132 41599 17184 41608
rect 17132 41565 17141 41599
rect 17141 41565 17175 41599
rect 17175 41565 17184 41599
rect 17132 41556 17184 41565
rect 20168 41599 20220 41608
rect 20168 41565 20177 41599
rect 20177 41565 20211 41599
rect 20211 41565 20220 41599
rect 20168 41556 20220 41565
rect 20628 41599 20680 41608
rect 20628 41565 20637 41599
rect 20637 41565 20671 41599
rect 20671 41565 20680 41599
rect 20628 41556 20680 41565
rect 20812 41599 20864 41608
rect 20812 41565 20821 41599
rect 20821 41565 20855 41599
rect 20855 41565 20864 41599
rect 20812 41556 20864 41565
rect 22836 41599 22888 41608
rect 22836 41565 22845 41599
rect 22845 41565 22879 41599
rect 22879 41565 22888 41599
rect 22836 41556 22888 41565
rect 26516 41556 26568 41608
rect 26792 41599 26844 41608
rect 26792 41565 26801 41599
rect 26801 41565 26835 41599
rect 26835 41565 26844 41599
rect 26792 41556 26844 41565
rect 16672 41488 16724 41540
rect 20536 41531 20588 41540
rect 20536 41497 20545 41531
rect 20545 41497 20579 41531
rect 20579 41497 20588 41531
rect 20536 41488 20588 41497
rect 23480 41488 23532 41540
rect 17040 41420 17092 41472
rect 21088 41420 21140 41472
rect 24400 41420 24452 41472
rect 26700 41463 26752 41472
rect 26700 41429 26709 41463
rect 26709 41429 26743 41463
rect 26743 41429 26752 41463
rect 26700 41420 26752 41429
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 16672 41259 16724 41268
rect 16672 41225 16681 41259
rect 16681 41225 16715 41259
rect 16715 41225 16724 41259
rect 16672 41216 16724 41225
rect 23480 41259 23532 41268
rect 23480 41225 23489 41259
rect 23489 41225 23523 41259
rect 23523 41225 23532 41259
rect 23480 41216 23532 41225
rect 16580 41148 16632 41200
rect 19616 41148 19668 41200
rect 17040 41012 17092 41064
rect 17592 41080 17644 41132
rect 20168 41080 20220 41132
rect 23388 41123 23440 41132
rect 23388 41089 23397 41123
rect 23397 41089 23431 41123
rect 23431 41089 23440 41123
rect 23388 41080 23440 41089
rect 26700 41148 26752 41200
rect 24124 41123 24176 41132
rect 24124 41089 24133 41123
rect 24133 41089 24167 41123
rect 24167 41089 24176 41123
rect 24124 41080 24176 41089
rect 26424 41123 26476 41132
rect 26424 41089 26433 41123
rect 26433 41089 26467 41123
rect 26467 41089 26476 41123
rect 26424 41080 26476 41089
rect 23204 41012 23256 41064
rect 21180 40944 21232 40996
rect 24584 41012 24636 41064
rect 26148 41012 26200 41064
rect 26976 41055 27028 41064
rect 26976 41021 26985 41055
rect 26985 41021 27019 41055
rect 27019 41021 27028 41055
rect 26976 41012 27028 41021
rect 17592 40876 17644 40928
rect 27160 40876 27212 40928
rect 27712 40876 27764 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 20536 40672 20588 40724
rect 21088 40715 21140 40724
rect 21088 40681 21097 40715
rect 21097 40681 21131 40715
rect 21131 40681 21140 40715
rect 21088 40672 21140 40681
rect 23204 40715 23256 40724
rect 23204 40681 23213 40715
rect 23213 40681 23247 40715
rect 23247 40681 23256 40715
rect 23204 40672 23256 40681
rect 20628 40604 20680 40656
rect 21180 40604 21232 40656
rect 17592 40468 17644 40520
rect 21088 40536 21140 40588
rect 20996 40511 21048 40520
rect 20996 40477 21005 40511
rect 21005 40477 21039 40511
rect 21039 40477 21048 40511
rect 20996 40468 21048 40477
rect 23480 40536 23532 40588
rect 24216 40672 24268 40724
rect 26608 40672 26660 40724
rect 26792 40672 26844 40724
rect 24124 40468 24176 40520
rect 24400 40511 24452 40520
rect 24400 40477 24409 40511
rect 24409 40477 24443 40511
rect 24443 40477 24452 40511
rect 24400 40468 24452 40477
rect 26332 40511 26384 40520
rect 26332 40477 26341 40511
rect 26341 40477 26375 40511
rect 26375 40477 26384 40511
rect 26332 40468 26384 40477
rect 26700 40536 26752 40588
rect 27160 40579 27212 40588
rect 27160 40545 27169 40579
rect 27169 40545 27203 40579
rect 27203 40545 27212 40579
rect 27160 40536 27212 40545
rect 27344 40579 27396 40588
rect 27344 40545 27353 40579
rect 27353 40545 27387 40579
rect 27387 40545 27396 40579
rect 27344 40536 27396 40545
rect 27436 40468 27488 40520
rect 26240 40400 26292 40452
rect 23940 40332 23992 40384
rect 24308 40332 24360 40384
rect 27252 40332 27304 40384
rect 27528 40375 27580 40384
rect 27528 40341 27537 40375
rect 27537 40341 27571 40375
rect 27571 40341 27580 40375
rect 27528 40332 27580 40341
rect 27896 40375 27948 40384
rect 27896 40341 27905 40375
rect 27905 40341 27939 40375
rect 27939 40341 27948 40375
rect 27896 40332 27948 40341
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 20996 40128 21048 40180
rect 23480 40128 23532 40180
rect 26148 40128 26200 40180
rect 26424 40128 26476 40180
rect 27896 40171 27948 40180
rect 27896 40137 27905 40171
rect 27905 40137 27939 40171
rect 27939 40137 27948 40171
rect 27896 40128 27948 40137
rect 9588 40060 9640 40112
rect 11060 39992 11112 40044
rect 12072 40035 12124 40044
rect 12072 40001 12081 40035
rect 12081 40001 12115 40035
rect 12115 40001 12124 40035
rect 12072 39992 12124 40001
rect 12624 39992 12676 40044
rect 19892 39992 19944 40044
rect 20076 39992 20128 40044
rect 9312 39967 9364 39976
rect 9312 39933 9321 39967
rect 9321 39933 9355 39967
rect 9355 39933 9364 39967
rect 9312 39924 9364 39933
rect 20168 39856 20220 39908
rect 20812 40035 20864 40044
rect 20812 40001 20821 40035
rect 20821 40001 20855 40035
rect 20855 40001 20864 40035
rect 20812 39992 20864 40001
rect 20996 40035 21048 40044
rect 20996 40001 21005 40035
rect 21005 40001 21039 40035
rect 21039 40001 21048 40035
rect 20996 39992 21048 40001
rect 21364 39992 21416 40044
rect 23112 39992 23164 40044
rect 21272 39856 21324 39908
rect 21640 39856 21692 39908
rect 23296 40035 23348 40044
rect 23296 40001 23305 40035
rect 23305 40001 23339 40035
rect 23339 40001 23348 40035
rect 23296 39992 23348 40001
rect 23940 40035 23992 40044
rect 23940 40001 23949 40035
rect 23949 40001 23983 40035
rect 23983 40001 23992 40035
rect 23940 39992 23992 40001
rect 27436 40103 27488 40112
rect 27436 40069 27445 40103
rect 27445 40069 27479 40103
rect 27479 40069 27488 40103
rect 27436 40060 27488 40069
rect 27712 40103 27764 40112
rect 27712 40069 27721 40103
rect 27721 40069 27755 40103
rect 27755 40069 27764 40103
rect 27712 40060 27764 40069
rect 24400 40035 24452 40044
rect 24400 40001 24409 40035
rect 24409 40001 24443 40035
rect 24443 40001 24452 40035
rect 24400 39992 24452 40001
rect 24676 40035 24728 40044
rect 24676 40001 24685 40035
rect 24685 40001 24719 40035
rect 24719 40001 24728 40035
rect 24676 39992 24728 40001
rect 26240 39992 26292 40044
rect 26700 39992 26752 40044
rect 23664 39967 23716 39976
rect 23664 39933 23673 39967
rect 23673 39933 23707 39967
rect 23707 39933 23716 39967
rect 23664 39924 23716 39933
rect 27896 39856 27948 39908
rect 8484 39788 8536 39840
rect 13452 39831 13504 39840
rect 13452 39797 13461 39831
rect 13461 39797 13495 39831
rect 13495 39797 13504 39831
rect 13452 39788 13504 39797
rect 19800 39788 19852 39840
rect 20444 39831 20496 39840
rect 20444 39797 20453 39831
rect 20453 39797 20487 39831
rect 20487 39797 20496 39831
rect 20444 39788 20496 39797
rect 20628 39788 20680 39840
rect 21364 39788 21416 39840
rect 24032 39788 24084 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 11060 39584 11112 39636
rect 17408 39584 17460 39636
rect 17592 39627 17644 39636
rect 17592 39593 17601 39627
rect 17601 39593 17635 39627
rect 17635 39593 17644 39627
rect 17592 39584 17644 39593
rect 18328 39584 18380 39636
rect 20168 39584 20220 39636
rect 20996 39584 21048 39636
rect 21088 39627 21140 39636
rect 21088 39593 21097 39627
rect 21097 39593 21131 39627
rect 21131 39593 21140 39627
rect 21088 39584 21140 39593
rect 21272 39584 21324 39636
rect 23572 39584 23624 39636
rect 23664 39584 23716 39636
rect 12072 39448 12124 39500
rect 16764 39491 16816 39500
rect 16764 39457 16773 39491
rect 16773 39457 16807 39491
rect 16807 39457 16816 39491
rect 16764 39448 16816 39457
rect 8484 39423 8536 39432
rect 8484 39389 8493 39423
rect 8493 39389 8527 39423
rect 8527 39389 8536 39423
rect 8484 39380 8536 39389
rect 8944 39423 8996 39432
rect 8944 39389 8953 39423
rect 8953 39389 8987 39423
rect 8987 39389 8996 39423
rect 8944 39380 8996 39389
rect 9588 39380 9640 39432
rect 12440 39380 12492 39432
rect 13360 39380 13412 39432
rect 17040 39448 17092 39500
rect 12256 39355 12308 39364
rect 12256 39321 12265 39355
rect 12265 39321 12299 39355
rect 12299 39321 12308 39355
rect 12256 39312 12308 39321
rect 13176 39312 13228 39364
rect 16212 39312 16264 39364
rect 17776 39312 17828 39364
rect 19800 39423 19852 39432
rect 19800 39389 19809 39423
rect 19809 39389 19843 39423
rect 19843 39389 19852 39423
rect 19800 39380 19852 39389
rect 19892 39423 19944 39432
rect 19892 39389 19901 39423
rect 19901 39389 19935 39423
rect 19935 39389 19944 39423
rect 19892 39380 19944 39389
rect 20076 39423 20128 39432
rect 20076 39389 20085 39423
rect 20085 39389 20119 39423
rect 20119 39389 20128 39423
rect 20076 39380 20128 39389
rect 20444 39491 20496 39500
rect 20444 39457 20453 39491
rect 20453 39457 20487 39491
rect 20487 39457 20496 39491
rect 20444 39448 20496 39457
rect 21272 39491 21324 39500
rect 21272 39457 21281 39491
rect 21281 39457 21315 39491
rect 21315 39457 21324 39491
rect 21272 39448 21324 39457
rect 24676 39516 24728 39568
rect 21364 39423 21416 39432
rect 21364 39389 21373 39423
rect 21373 39389 21407 39423
rect 21407 39389 21416 39423
rect 21364 39380 21416 39389
rect 21640 39423 21692 39432
rect 21640 39389 21649 39423
rect 21649 39389 21683 39423
rect 21683 39389 21692 39423
rect 21640 39380 21692 39389
rect 9680 39244 9732 39296
rect 10324 39287 10376 39296
rect 10324 39253 10333 39287
rect 10333 39253 10367 39287
rect 10367 39253 10376 39287
rect 10324 39244 10376 39253
rect 14556 39244 14608 39296
rect 17224 39287 17276 39296
rect 17224 39253 17233 39287
rect 17233 39253 17267 39287
rect 17267 39253 17276 39287
rect 17224 39244 17276 39253
rect 18512 39244 18564 39296
rect 19432 39287 19484 39296
rect 19432 39253 19441 39287
rect 19441 39253 19475 39287
rect 19475 39253 19484 39287
rect 19432 39244 19484 39253
rect 23572 39355 23624 39364
rect 23572 39321 23581 39355
rect 23581 39321 23615 39355
rect 23615 39321 23624 39355
rect 24032 39423 24084 39432
rect 24032 39389 24041 39423
rect 24041 39389 24075 39423
rect 24075 39389 24084 39423
rect 24032 39380 24084 39389
rect 24216 39423 24268 39432
rect 24216 39389 24225 39423
rect 24225 39389 24259 39423
rect 24259 39389 24268 39423
rect 24216 39380 24268 39389
rect 23572 39312 23624 39321
rect 23112 39244 23164 39296
rect 23296 39244 23348 39296
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 9312 39040 9364 39092
rect 13176 39083 13228 39092
rect 13176 39049 13185 39083
rect 13185 39049 13219 39083
rect 13219 39049 13228 39083
rect 13176 39040 13228 39049
rect 16212 39083 16264 39092
rect 16212 39049 16221 39083
rect 16221 39049 16255 39083
rect 16255 39049 16264 39083
rect 16212 39040 16264 39049
rect 8944 38972 8996 39024
rect 7932 38947 7984 38956
rect 7932 38913 7966 38947
rect 7966 38913 7984 38947
rect 7932 38904 7984 38913
rect 9588 38947 9640 38956
rect 9588 38913 9597 38947
rect 9597 38913 9631 38947
rect 9631 38913 9640 38947
rect 9588 38904 9640 38913
rect 9864 38947 9916 38956
rect 9864 38913 9898 38947
rect 9898 38913 9916 38947
rect 9864 38904 9916 38913
rect 13360 38947 13412 38956
rect 13360 38913 13369 38947
rect 13369 38913 13403 38947
rect 13403 38913 13412 38947
rect 13360 38904 13412 38913
rect 13452 38947 13504 38956
rect 13452 38913 13461 38947
rect 13461 38913 13495 38947
rect 13495 38913 13504 38947
rect 13452 38904 13504 38913
rect 14556 38947 14608 38956
rect 14556 38913 14565 38947
rect 14565 38913 14599 38947
rect 14599 38913 14608 38947
rect 14556 38904 14608 38913
rect 14280 38836 14332 38888
rect 16028 38947 16080 38956
rect 16028 38913 16037 38947
rect 16037 38913 16071 38947
rect 16071 38913 16080 38947
rect 16028 38904 16080 38913
rect 16212 38947 16264 38956
rect 16212 38913 16221 38947
rect 16221 38913 16255 38947
rect 16255 38913 16264 38947
rect 16212 38904 16264 38913
rect 16856 39040 16908 39092
rect 17132 38972 17184 39024
rect 10600 38700 10652 38752
rect 15384 38700 15436 38752
rect 18328 38947 18380 38956
rect 18328 38913 18337 38947
rect 18337 38913 18371 38947
rect 18371 38913 18380 38947
rect 18328 38904 18380 38913
rect 18604 38947 18656 38956
rect 18604 38913 18613 38947
rect 18613 38913 18647 38947
rect 18647 38913 18656 38947
rect 18604 38904 18656 38913
rect 18236 38768 18288 38820
rect 18880 38879 18932 38888
rect 18880 38845 18889 38879
rect 18889 38845 18923 38879
rect 18923 38845 18932 38879
rect 18880 38836 18932 38845
rect 19432 39040 19484 39092
rect 19524 38972 19576 39024
rect 19892 38904 19944 38956
rect 20260 38904 20312 38956
rect 23296 38904 23348 38956
rect 16580 38700 16632 38752
rect 16672 38700 16724 38752
rect 17776 38700 17828 38752
rect 18144 38743 18196 38752
rect 18144 38709 18153 38743
rect 18153 38709 18187 38743
rect 18187 38709 18196 38743
rect 18144 38700 18196 38709
rect 18696 38743 18748 38752
rect 18696 38709 18705 38743
rect 18705 38709 18739 38743
rect 18739 38709 18748 38743
rect 18696 38700 18748 38709
rect 21180 38879 21232 38888
rect 21180 38845 21189 38879
rect 21189 38845 21223 38879
rect 21223 38845 21232 38879
rect 21180 38836 21232 38845
rect 23112 38879 23164 38888
rect 23112 38845 23121 38879
rect 23121 38845 23155 38879
rect 23155 38845 23164 38879
rect 23112 38836 23164 38845
rect 20444 38811 20496 38820
rect 20444 38777 20453 38811
rect 20453 38777 20487 38811
rect 20487 38777 20496 38811
rect 20444 38768 20496 38777
rect 20812 38768 20864 38820
rect 23572 38811 23624 38820
rect 23572 38777 23581 38811
rect 23581 38777 23615 38811
rect 23615 38777 23624 38811
rect 23572 38768 23624 38777
rect 19340 38700 19392 38752
rect 20536 38743 20588 38752
rect 20536 38709 20545 38743
rect 20545 38709 20579 38743
rect 20579 38709 20588 38743
rect 20536 38700 20588 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 7932 38496 7984 38548
rect 9864 38539 9916 38548
rect 9864 38505 9873 38539
rect 9873 38505 9907 38539
rect 9907 38505 9916 38539
rect 9864 38496 9916 38505
rect 14280 38539 14332 38548
rect 14280 38505 14289 38539
rect 14289 38505 14323 38539
rect 14323 38505 14332 38539
rect 14280 38496 14332 38505
rect 16672 38496 16724 38548
rect 16764 38539 16816 38548
rect 16764 38505 16773 38539
rect 16773 38505 16807 38539
rect 16807 38505 16816 38539
rect 16764 38496 16816 38505
rect 16856 38539 16908 38548
rect 16856 38505 16865 38539
rect 16865 38505 16899 38539
rect 16899 38505 16908 38539
rect 16856 38496 16908 38505
rect 19524 38539 19576 38548
rect 19524 38505 19533 38539
rect 19533 38505 19567 38539
rect 19567 38505 19576 38539
rect 19524 38496 19576 38505
rect 20076 38539 20128 38548
rect 20076 38505 20085 38539
rect 20085 38505 20119 38539
rect 20119 38505 20128 38539
rect 20076 38496 20128 38505
rect 26884 38496 26936 38548
rect 27344 38496 27396 38548
rect 13452 38403 13504 38412
rect 13452 38369 13461 38403
rect 13461 38369 13495 38403
rect 13495 38369 13504 38403
rect 13452 38360 13504 38369
rect 16028 38428 16080 38480
rect 8300 38335 8352 38344
rect 8300 38301 8309 38335
rect 8309 38301 8343 38335
rect 8343 38301 8352 38335
rect 8300 38292 8352 38301
rect 8576 38292 8628 38344
rect 9680 38335 9732 38344
rect 9680 38301 9689 38335
rect 9689 38301 9723 38335
rect 9723 38301 9732 38335
rect 9680 38292 9732 38301
rect 10600 38335 10652 38344
rect 10600 38301 10609 38335
rect 10609 38301 10643 38335
rect 10643 38301 10652 38335
rect 10600 38292 10652 38301
rect 10324 38224 10376 38276
rect 12532 38292 12584 38344
rect 13728 38292 13780 38344
rect 14556 38335 14608 38344
rect 14556 38301 14565 38335
rect 14565 38301 14599 38335
rect 14599 38301 14608 38335
rect 14556 38292 14608 38301
rect 14648 38335 14700 38344
rect 14648 38301 14657 38335
rect 14657 38301 14691 38335
rect 14691 38301 14700 38335
rect 14648 38292 14700 38301
rect 15384 38335 15436 38344
rect 15384 38301 15393 38335
rect 15393 38301 15427 38335
rect 15427 38301 15436 38335
rect 15384 38292 15436 38301
rect 18144 38428 18196 38480
rect 17224 38360 17276 38412
rect 17408 38403 17460 38412
rect 17408 38369 17417 38403
rect 17417 38369 17451 38403
rect 17451 38369 17460 38403
rect 17408 38360 17460 38369
rect 16948 38292 17000 38344
rect 18696 38360 18748 38412
rect 17684 38335 17736 38344
rect 17684 38301 17693 38335
rect 17693 38301 17727 38335
rect 17727 38301 17736 38335
rect 17684 38292 17736 38301
rect 10140 38156 10192 38208
rect 14280 38156 14332 38208
rect 16212 38156 16264 38208
rect 16488 38156 16540 38208
rect 18236 38335 18288 38344
rect 18236 38301 18245 38335
rect 18245 38301 18279 38335
rect 18279 38301 18288 38335
rect 18236 38292 18288 38301
rect 20536 38428 20588 38480
rect 20628 38360 20680 38412
rect 27160 38403 27212 38412
rect 27160 38369 27169 38403
rect 27169 38369 27203 38403
rect 27203 38369 27212 38403
rect 27160 38360 27212 38369
rect 18880 38224 18932 38276
rect 19616 38224 19668 38276
rect 20444 38292 20496 38344
rect 27528 38292 27580 38344
rect 18328 38199 18380 38208
rect 18328 38165 18337 38199
rect 18337 38165 18371 38199
rect 18371 38165 18380 38199
rect 18328 38156 18380 38165
rect 20260 38156 20312 38208
rect 27068 38156 27120 38208
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 8576 37995 8628 38004
rect 8576 37961 8585 37995
rect 8585 37961 8619 37995
rect 8619 37961 8628 37995
rect 8576 37952 8628 37961
rect 10600 37952 10652 38004
rect 16028 37952 16080 38004
rect 17684 37952 17736 38004
rect 17776 37952 17828 38004
rect 9312 37884 9364 37936
rect 10324 37884 10376 37936
rect 12440 37927 12492 37936
rect 12440 37893 12449 37927
rect 12449 37893 12483 37927
rect 12483 37893 12492 37927
rect 12440 37884 12492 37893
rect 12624 37884 12676 37936
rect 9680 37859 9732 37868
rect 9680 37825 9689 37859
rect 9689 37825 9723 37859
rect 9723 37825 9732 37859
rect 9680 37816 9732 37825
rect 8484 37748 8536 37800
rect 13268 37816 13320 37868
rect 13728 37816 13780 37868
rect 14556 37884 14608 37936
rect 18328 37884 18380 37936
rect 19616 37952 19668 38004
rect 20536 37952 20588 38004
rect 23572 37952 23624 38004
rect 27160 37952 27212 38004
rect 14280 37859 14332 37868
rect 14280 37825 14289 37859
rect 14289 37825 14323 37859
rect 14323 37825 14332 37859
rect 14280 37816 14332 37825
rect 11152 37791 11204 37800
rect 11152 37757 11161 37791
rect 11161 37757 11195 37791
rect 11195 37757 11204 37791
rect 11152 37748 11204 37757
rect 12716 37748 12768 37800
rect 13452 37748 13504 37800
rect 14648 37816 14700 37868
rect 23664 37859 23716 37868
rect 23664 37825 23673 37859
rect 23673 37825 23707 37859
rect 23707 37825 23716 37859
rect 23664 37816 23716 37825
rect 27160 37816 27212 37868
rect 27344 37859 27396 37868
rect 27344 37825 27353 37859
rect 27353 37825 27387 37859
rect 27387 37825 27396 37859
rect 27344 37816 27396 37825
rect 16488 37748 16540 37800
rect 26240 37748 26292 37800
rect 9772 37612 9824 37664
rect 10508 37612 10560 37664
rect 16948 37655 17000 37664
rect 16948 37621 16957 37655
rect 16957 37621 16991 37655
rect 16991 37621 17000 37655
rect 16948 37612 17000 37621
rect 24584 37680 24636 37732
rect 26884 37680 26936 37732
rect 23296 37655 23348 37664
rect 23296 37621 23305 37655
rect 23305 37621 23339 37655
rect 23339 37621 23348 37655
rect 23296 37612 23348 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 8300 37408 8352 37460
rect 10140 37451 10192 37460
rect 10140 37417 10149 37451
rect 10149 37417 10183 37451
rect 10183 37417 10192 37451
rect 10140 37408 10192 37417
rect 23756 37408 23808 37460
rect 9680 37340 9732 37392
rect 8392 37204 8444 37256
rect 9312 37272 9364 37324
rect 10324 37315 10376 37324
rect 10324 37281 10333 37315
rect 10333 37281 10367 37315
rect 10367 37281 10376 37315
rect 10324 37272 10376 37281
rect 8024 37136 8076 37188
rect 9220 37247 9272 37256
rect 9220 37213 9229 37247
rect 9229 37213 9263 37247
rect 9263 37213 9272 37247
rect 9220 37204 9272 37213
rect 9680 37204 9732 37256
rect 22836 37247 22888 37256
rect 22836 37213 22845 37247
rect 22845 37213 22879 37247
rect 22879 37213 22888 37247
rect 22836 37204 22888 37213
rect 9312 37136 9364 37188
rect 10968 37179 11020 37188
rect 10968 37145 11002 37179
rect 11002 37145 11020 37179
rect 10968 37136 11020 37145
rect 11060 37136 11112 37188
rect 12440 37179 12492 37188
rect 12440 37145 12474 37179
rect 12474 37145 12492 37179
rect 12440 37136 12492 37145
rect 23204 37136 23256 37188
rect 24400 37247 24452 37256
rect 24400 37213 24409 37247
rect 24409 37213 24443 37247
rect 24443 37213 24452 37247
rect 24400 37204 24452 37213
rect 26516 37204 26568 37256
rect 26884 37247 26936 37256
rect 26884 37213 26893 37247
rect 26893 37213 26927 37247
rect 26927 37213 26936 37247
rect 26884 37204 26936 37213
rect 27068 37247 27120 37256
rect 27068 37213 27077 37247
rect 27077 37213 27111 37247
rect 27111 37213 27120 37247
rect 27068 37204 27120 37213
rect 27160 37247 27212 37256
rect 27160 37213 27169 37247
rect 27169 37213 27203 37247
rect 27203 37213 27212 37247
rect 27160 37204 27212 37213
rect 28448 37247 28500 37256
rect 28448 37213 28457 37247
rect 28457 37213 28491 37247
rect 28491 37213 28500 37247
rect 28448 37204 28500 37213
rect 11152 37068 11204 37120
rect 12532 37068 12584 37120
rect 14280 37068 14332 37120
rect 24032 37068 24084 37120
rect 24400 37068 24452 37120
rect 26608 37179 26660 37188
rect 26608 37145 26617 37179
rect 26617 37145 26651 37179
rect 26651 37145 26660 37179
rect 26608 37136 26660 37145
rect 26884 37068 26936 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 8024 36907 8076 36916
rect 8024 36873 8033 36907
rect 8033 36873 8067 36907
rect 8067 36873 8076 36907
rect 8024 36864 8076 36873
rect 8484 36728 8536 36780
rect 9312 36660 9364 36712
rect 10968 36864 11020 36916
rect 10508 36839 10560 36848
rect 10508 36805 10517 36839
rect 10517 36805 10551 36839
rect 10551 36805 10560 36839
rect 10508 36796 10560 36805
rect 11796 36796 11848 36848
rect 9772 36728 9824 36780
rect 9680 36703 9732 36712
rect 9680 36669 9689 36703
rect 9689 36669 9723 36703
rect 9723 36669 9732 36703
rect 9680 36660 9732 36669
rect 8300 36592 8352 36644
rect 12440 36864 12492 36916
rect 23204 36907 23256 36916
rect 23204 36873 23213 36907
rect 23213 36873 23247 36907
rect 23247 36873 23256 36907
rect 23204 36864 23256 36873
rect 27344 36864 27396 36916
rect 12624 36796 12676 36848
rect 12532 36771 12584 36780
rect 12532 36737 12541 36771
rect 12541 36737 12575 36771
rect 12575 36737 12584 36771
rect 12532 36728 12584 36737
rect 19340 36728 19392 36780
rect 22836 36728 22888 36780
rect 23388 36796 23440 36848
rect 26608 36796 26660 36848
rect 23296 36771 23348 36780
rect 23296 36737 23305 36771
rect 23305 36737 23339 36771
rect 23339 36737 23348 36771
rect 23296 36728 23348 36737
rect 26976 36771 27028 36780
rect 26976 36737 26985 36771
rect 26985 36737 27019 36771
rect 27019 36737 27028 36771
rect 26976 36728 27028 36737
rect 28448 36524 28500 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 9220 36184 9272 36236
rect 9496 36227 9548 36236
rect 9496 36193 9505 36227
rect 9505 36193 9539 36227
rect 9539 36193 9548 36227
rect 9496 36184 9548 36193
rect 22836 36184 22888 36236
rect 12256 36048 12308 36100
rect 19892 36048 19944 36100
rect 8944 36023 8996 36032
rect 8944 35989 8953 36023
rect 8953 35989 8987 36023
rect 8987 35989 8996 36023
rect 8944 35980 8996 35989
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 6920 35776 6972 35828
rect 8392 35708 8444 35760
rect 6368 35615 6420 35624
rect 6368 35581 6377 35615
rect 6377 35581 6411 35615
rect 6411 35581 6420 35615
rect 6368 35572 6420 35581
rect 8944 35683 8996 35692
rect 8944 35649 8953 35683
rect 8953 35649 8987 35683
rect 8987 35649 8996 35683
rect 8944 35640 8996 35649
rect 9312 35819 9364 35828
rect 9312 35785 9321 35819
rect 9321 35785 9355 35819
rect 9355 35785 9364 35819
rect 9312 35776 9364 35785
rect 9680 35708 9732 35760
rect 12072 35708 12124 35760
rect 18604 35708 18656 35760
rect 11888 35640 11940 35692
rect 18880 35640 18932 35692
rect 20352 35640 20404 35692
rect 28264 35683 28316 35692
rect 28264 35649 28273 35683
rect 28273 35649 28307 35683
rect 28307 35649 28316 35683
rect 28264 35640 28316 35649
rect 10692 35615 10744 35624
rect 10692 35581 10701 35615
rect 10701 35581 10735 35615
rect 10735 35581 10744 35615
rect 10692 35572 10744 35581
rect 26792 35572 26844 35624
rect 9496 35504 9548 35556
rect 20720 35436 20772 35488
rect 27620 35479 27672 35488
rect 27620 35445 27629 35479
rect 27629 35445 27663 35479
rect 27663 35445 27672 35479
rect 27620 35436 27672 35445
rect 28448 35479 28500 35488
rect 28448 35445 28457 35479
rect 28457 35445 28491 35479
rect 28491 35445 28500 35479
rect 28448 35436 28500 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 6368 35275 6420 35284
rect 6368 35241 6377 35275
rect 6377 35241 6411 35275
rect 6411 35241 6420 35275
rect 6368 35232 6420 35241
rect 11796 35275 11848 35284
rect 11796 35241 11805 35275
rect 11805 35241 11839 35275
rect 11839 35241 11848 35275
rect 11796 35232 11848 35241
rect 11888 35275 11940 35284
rect 11888 35241 11897 35275
rect 11897 35241 11931 35275
rect 11931 35241 11940 35275
rect 11888 35232 11940 35241
rect 28264 35275 28316 35284
rect 28264 35241 28273 35275
rect 28273 35241 28307 35275
rect 28307 35241 28316 35275
rect 28264 35232 28316 35241
rect 7012 35139 7064 35148
rect 7012 35105 7021 35139
rect 7021 35105 7055 35139
rect 7055 35105 7064 35139
rect 7012 35096 7064 35105
rect 8300 35096 8352 35148
rect 18880 35164 18932 35216
rect 19524 35139 19576 35148
rect 19524 35105 19533 35139
rect 19533 35105 19567 35139
rect 19567 35105 19576 35139
rect 19524 35096 19576 35105
rect 11152 35071 11204 35080
rect 11152 35037 11161 35071
rect 11161 35037 11195 35071
rect 11195 35037 11204 35071
rect 11152 35028 11204 35037
rect 12072 35071 12124 35080
rect 12072 35037 12081 35071
rect 12081 35037 12115 35071
rect 12115 35037 12124 35071
rect 12072 35028 12124 35037
rect 19432 35071 19484 35080
rect 19432 35037 19441 35071
rect 19441 35037 19475 35071
rect 19475 35037 19484 35071
rect 19432 35028 19484 35037
rect 8392 35003 8444 35012
rect 8392 34969 8401 35003
rect 8401 34969 8435 35003
rect 8435 34969 8444 35003
rect 8392 34960 8444 34969
rect 12164 34960 12216 35012
rect 18328 34960 18380 35012
rect 20812 35028 20864 35080
rect 20904 35071 20956 35080
rect 20904 35037 20913 35071
rect 20913 35037 20947 35071
rect 20947 35037 20956 35071
rect 20904 35028 20956 35037
rect 26976 35028 27028 35080
rect 27620 35028 27672 35080
rect 22008 34960 22060 35012
rect 8852 34892 8904 34944
rect 10692 34892 10744 34944
rect 19340 34892 19392 34944
rect 20628 34892 20680 34944
rect 20996 34892 21048 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 7012 34688 7064 34740
rect 11152 34688 11204 34740
rect 20352 34731 20404 34740
rect 20352 34697 20361 34731
rect 20361 34697 20395 34731
rect 20395 34697 20404 34731
rect 20352 34688 20404 34697
rect 20812 34688 20864 34740
rect 25228 34688 25280 34740
rect 27344 34688 27396 34740
rect 4620 34484 4672 34536
rect 9680 34620 9732 34672
rect 18328 34620 18380 34672
rect 16212 34595 16264 34604
rect 16212 34561 16230 34595
rect 16230 34561 16264 34595
rect 16212 34552 16264 34561
rect 18512 34595 18564 34604
rect 18512 34561 18521 34595
rect 18521 34561 18555 34595
rect 18555 34561 18564 34595
rect 18512 34552 18564 34561
rect 18604 34595 18656 34604
rect 18604 34561 18613 34595
rect 18613 34561 18647 34595
rect 18647 34561 18656 34595
rect 18604 34552 18656 34561
rect 21364 34663 21416 34672
rect 21364 34629 21373 34663
rect 21373 34629 21407 34663
rect 21407 34629 21416 34663
rect 21364 34620 21416 34629
rect 18880 34595 18932 34604
rect 18880 34561 18889 34595
rect 18889 34561 18923 34595
rect 18923 34561 18932 34595
rect 18880 34552 18932 34561
rect 19432 34552 19484 34604
rect 20260 34552 20312 34604
rect 8852 34484 8904 34536
rect 17776 34484 17828 34536
rect 19340 34416 19392 34468
rect 19616 34527 19668 34536
rect 19616 34493 19625 34527
rect 19625 34493 19659 34527
rect 19659 34493 19668 34527
rect 19616 34484 19668 34493
rect 15016 34348 15068 34400
rect 19524 34348 19576 34400
rect 22008 34595 22060 34604
rect 22008 34561 22017 34595
rect 22017 34561 22051 34595
rect 22051 34561 22060 34595
rect 22008 34552 22060 34561
rect 22928 34620 22980 34672
rect 24308 34620 24360 34672
rect 26792 34663 26844 34672
rect 26792 34629 26801 34663
rect 26801 34629 26835 34663
rect 26835 34629 26844 34663
rect 26792 34620 26844 34629
rect 22100 34484 22152 34536
rect 23664 34552 23716 34604
rect 26516 34552 26568 34604
rect 26976 34595 27028 34604
rect 26976 34561 26985 34595
rect 26985 34561 27019 34595
rect 27019 34561 27028 34595
rect 26976 34552 27028 34561
rect 24860 34484 24912 34536
rect 25596 34484 25648 34536
rect 27436 34552 27488 34604
rect 27252 34527 27304 34536
rect 27252 34493 27261 34527
rect 27261 34493 27295 34527
rect 27295 34493 27304 34527
rect 27252 34484 27304 34493
rect 27988 34484 28040 34536
rect 22928 34416 22980 34468
rect 26608 34459 26660 34468
rect 26608 34425 26617 34459
rect 26617 34425 26651 34459
rect 26651 34425 26660 34459
rect 26608 34416 26660 34425
rect 25412 34348 25464 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 16212 34187 16264 34196
rect 16212 34153 16221 34187
rect 16221 34153 16255 34187
rect 16255 34153 16264 34187
rect 16212 34144 16264 34153
rect 17776 34144 17828 34196
rect 18696 34076 18748 34128
rect 15016 33940 15068 33992
rect 17500 34008 17552 34060
rect 15108 33872 15160 33924
rect 16672 33940 16724 33992
rect 18604 34008 18656 34060
rect 19156 34008 19208 34060
rect 18052 33915 18104 33924
rect 18052 33881 18061 33915
rect 18061 33881 18095 33915
rect 18095 33881 18104 33915
rect 18052 33872 18104 33881
rect 15936 33847 15988 33856
rect 15936 33813 15945 33847
rect 15945 33813 15979 33847
rect 15979 33813 15988 33847
rect 15936 33804 15988 33813
rect 17868 33847 17920 33856
rect 17868 33813 17877 33847
rect 17877 33813 17911 33847
rect 17911 33813 17920 33847
rect 17868 33804 17920 33813
rect 22100 34008 22152 34060
rect 23204 34144 23256 34196
rect 26976 34144 27028 34196
rect 27988 34051 28040 34060
rect 27988 34017 27997 34051
rect 27997 34017 28031 34051
rect 28031 34017 28040 34051
rect 27988 34008 28040 34017
rect 21180 33940 21232 33992
rect 21272 33940 21324 33992
rect 19984 33872 20036 33924
rect 22468 33872 22520 33924
rect 18880 33804 18932 33856
rect 19248 33847 19300 33856
rect 19248 33813 19257 33847
rect 19257 33813 19291 33847
rect 19291 33813 19300 33847
rect 19248 33804 19300 33813
rect 22284 33804 22336 33856
rect 25228 33983 25280 33992
rect 25228 33949 25237 33983
rect 25237 33949 25271 33983
rect 25271 33949 25280 33983
rect 25228 33940 25280 33949
rect 25412 33983 25464 33992
rect 25412 33949 25421 33983
rect 25421 33949 25455 33983
rect 25455 33949 25464 33983
rect 25412 33940 25464 33949
rect 25596 33983 25648 33992
rect 25596 33949 25605 33983
rect 25605 33949 25639 33983
rect 25639 33949 25648 33983
rect 25596 33940 25648 33949
rect 22928 33915 22980 33924
rect 22928 33881 22937 33915
rect 22937 33881 22971 33915
rect 22971 33881 22980 33915
rect 22928 33872 22980 33881
rect 27252 33872 27304 33924
rect 24032 33804 24084 33856
rect 26516 33804 26568 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 4620 33600 4672 33652
rect 15476 33532 15528 33584
rect 16672 33643 16724 33652
rect 16672 33609 16681 33643
rect 16681 33609 16715 33643
rect 16715 33609 16724 33643
rect 16672 33600 16724 33609
rect 17592 33643 17644 33652
rect 17592 33609 17601 33643
rect 17601 33609 17635 33643
rect 17635 33609 17644 33643
rect 17592 33600 17644 33609
rect 19156 33643 19208 33652
rect 19156 33609 19165 33643
rect 19165 33609 19199 33643
rect 19199 33609 19208 33643
rect 19156 33600 19208 33609
rect 3516 33507 3568 33516
rect 3516 33473 3525 33507
rect 3525 33473 3559 33507
rect 3559 33473 3568 33507
rect 3516 33464 3568 33473
rect 13268 33464 13320 33516
rect 15016 33507 15068 33516
rect 15016 33473 15025 33507
rect 15025 33473 15059 33507
rect 15059 33473 15068 33507
rect 15016 33464 15068 33473
rect 15108 33507 15160 33516
rect 15108 33473 15120 33507
rect 15120 33473 15154 33507
rect 15154 33473 15160 33507
rect 15108 33464 15160 33473
rect 17868 33532 17920 33584
rect 18144 33532 18196 33584
rect 21180 33643 21232 33652
rect 21180 33609 21189 33643
rect 21189 33609 21223 33643
rect 21223 33609 21232 33643
rect 21180 33600 21232 33609
rect 23204 33643 23256 33652
rect 23204 33609 23213 33643
rect 23213 33609 23247 33643
rect 23247 33609 23256 33643
rect 23204 33600 23256 33609
rect 2964 33396 3016 33448
rect 8852 33396 8904 33448
rect 13912 33371 13964 33380
rect 13912 33337 13921 33371
rect 13921 33337 13955 33371
rect 13955 33337 13964 33371
rect 15292 33396 15344 33448
rect 17500 33507 17552 33516
rect 17500 33473 17509 33507
rect 17509 33473 17543 33507
rect 17543 33473 17552 33507
rect 17500 33464 17552 33473
rect 17776 33507 17828 33516
rect 17776 33473 17785 33507
rect 17785 33473 17819 33507
rect 17819 33473 17828 33507
rect 17776 33464 17828 33473
rect 17224 33439 17276 33448
rect 17224 33405 17233 33439
rect 17233 33405 17267 33439
rect 17267 33405 17276 33439
rect 17224 33396 17276 33405
rect 19248 33464 19300 33516
rect 19892 33575 19944 33584
rect 19892 33541 19901 33575
rect 19901 33541 19935 33575
rect 19935 33541 19944 33575
rect 19892 33532 19944 33541
rect 22100 33507 22152 33516
rect 22100 33473 22134 33507
rect 22134 33473 22152 33507
rect 22100 33464 22152 33473
rect 22468 33464 22520 33516
rect 26608 33464 26660 33516
rect 20996 33396 21048 33448
rect 21180 33396 21232 33448
rect 13912 33328 13964 33337
rect 15384 33328 15436 33380
rect 15936 33328 15988 33380
rect 14004 33303 14056 33312
rect 14004 33269 14013 33303
rect 14013 33269 14047 33303
rect 14047 33269 14056 33303
rect 14004 33260 14056 33269
rect 19524 33260 19576 33312
rect 21272 33260 21324 33312
rect 23296 33303 23348 33312
rect 23296 33269 23305 33303
rect 23305 33269 23339 33303
rect 23339 33269 23348 33303
rect 23296 33260 23348 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 3516 33056 3568 33108
rect 13268 33099 13320 33108
rect 13268 33065 13277 33099
rect 13277 33065 13311 33099
rect 13311 33065 13320 33099
rect 13268 33056 13320 33065
rect 12532 32988 12584 33040
rect 13636 33056 13688 33108
rect 15108 33056 15160 33108
rect 19616 33056 19668 33108
rect 21272 33099 21324 33108
rect 21272 33065 21281 33099
rect 21281 33065 21315 33099
rect 21315 33065 21324 33099
rect 21272 33056 21324 33065
rect 22100 33056 22152 33108
rect 22928 33056 22980 33108
rect 14096 32988 14148 33040
rect 21180 32988 21232 33040
rect 12900 32963 12952 32972
rect 12900 32929 12909 32963
rect 12909 32929 12943 32963
rect 12943 32929 12952 32963
rect 12900 32920 12952 32929
rect 16580 32920 16632 32972
rect 17224 32920 17276 32972
rect 18604 32920 18656 32972
rect 21824 32963 21876 32972
rect 21824 32929 21833 32963
rect 21833 32929 21867 32963
rect 21867 32929 21876 32963
rect 21824 32920 21876 32929
rect 24860 33056 24912 33108
rect 848 32852 900 32904
rect 11888 32852 11940 32904
rect 12440 32895 12492 32904
rect 12440 32861 12449 32895
rect 12449 32861 12483 32895
rect 12483 32861 12492 32895
rect 12440 32852 12492 32861
rect 12624 32852 12676 32904
rect 14004 32852 14056 32904
rect 15292 32895 15344 32904
rect 15292 32861 15301 32895
rect 15301 32861 15335 32895
rect 15335 32861 15344 32895
rect 15292 32852 15344 32861
rect 15384 32895 15436 32904
rect 15384 32861 15393 32895
rect 15393 32861 15427 32895
rect 15427 32861 15436 32895
rect 15384 32852 15436 32861
rect 15476 32852 15528 32904
rect 18696 32895 18748 32904
rect 18696 32861 18705 32895
rect 18705 32861 18739 32895
rect 18739 32861 18748 32895
rect 18696 32852 18748 32861
rect 14188 32784 14240 32836
rect 20720 32827 20772 32836
rect 20720 32793 20738 32827
rect 20738 32793 20772 32827
rect 20720 32784 20772 32793
rect 13820 32716 13872 32768
rect 15568 32716 15620 32768
rect 19248 32716 19300 32768
rect 19524 32716 19576 32768
rect 23296 32852 23348 32904
rect 24032 32895 24084 32904
rect 24032 32861 24041 32895
rect 24041 32861 24075 32895
rect 24075 32861 24084 32895
rect 24032 32852 24084 32861
rect 24308 32852 24360 32904
rect 24860 32963 24912 32972
rect 24860 32929 24869 32963
rect 24869 32929 24903 32963
rect 24903 32929 24912 32963
rect 24860 32920 24912 32929
rect 22192 32784 22244 32836
rect 22376 32784 22428 32836
rect 22284 32716 22336 32768
rect 23296 32759 23348 32768
rect 23296 32725 23305 32759
rect 23305 32725 23339 32759
rect 23339 32725 23348 32759
rect 23296 32716 23348 32725
rect 24216 32716 24268 32768
rect 26148 32852 26200 32904
rect 27988 32920 28040 32972
rect 26792 32852 26844 32904
rect 25596 32784 25648 32836
rect 25688 32784 25740 32836
rect 24768 32716 24820 32768
rect 26792 32759 26844 32768
rect 26792 32725 26794 32759
rect 26794 32725 26828 32759
rect 26828 32725 26844 32759
rect 26792 32716 26844 32725
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 12900 32512 12952 32564
rect 15292 32512 15344 32564
rect 19984 32512 20036 32564
rect 20720 32555 20772 32564
rect 20720 32521 20729 32555
rect 20729 32521 20763 32555
rect 20763 32521 20772 32555
rect 20720 32512 20772 32521
rect 22192 32555 22244 32564
rect 22192 32521 22201 32555
rect 22201 32521 22235 32555
rect 22235 32521 22244 32555
rect 22192 32512 22244 32521
rect 24860 32512 24912 32564
rect 25596 32512 25648 32564
rect 26056 32512 26108 32564
rect 27988 32512 28040 32564
rect 13820 32444 13872 32496
rect 12808 32376 12860 32428
rect 13636 32376 13688 32428
rect 12532 32308 12584 32360
rect 13084 32351 13136 32360
rect 13084 32317 13093 32351
rect 13093 32317 13127 32351
rect 13127 32317 13136 32351
rect 13084 32308 13136 32317
rect 13176 32351 13228 32360
rect 13176 32317 13185 32351
rect 13185 32317 13219 32351
rect 13219 32317 13228 32351
rect 13176 32308 13228 32317
rect 13912 32376 13964 32428
rect 14096 32419 14148 32428
rect 14096 32385 14105 32419
rect 14105 32385 14139 32419
rect 14139 32385 14148 32419
rect 14096 32376 14148 32385
rect 14188 32419 14240 32428
rect 14188 32385 14197 32419
rect 14197 32385 14231 32419
rect 14231 32385 14240 32419
rect 14188 32376 14240 32385
rect 19248 32419 19300 32428
rect 19248 32385 19257 32419
rect 19257 32385 19291 32419
rect 19291 32385 19300 32419
rect 19248 32376 19300 32385
rect 21272 32444 21324 32496
rect 21824 32444 21876 32496
rect 20812 32419 20864 32428
rect 20812 32385 20821 32419
rect 20821 32385 20855 32419
rect 20855 32385 20864 32419
rect 20812 32376 20864 32385
rect 20996 32419 21048 32428
rect 20996 32385 21005 32419
rect 21005 32385 21039 32419
rect 21039 32385 21048 32419
rect 20996 32376 21048 32385
rect 22376 32419 22428 32428
rect 22376 32385 22385 32419
rect 22385 32385 22419 32419
rect 22419 32385 22428 32419
rect 22376 32376 22428 32385
rect 22468 32376 22520 32428
rect 23296 32376 23348 32428
rect 24400 32376 24452 32428
rect 25412 32419 25464 32428
rect 25412 32385 25446 32419
rect 25446 32385 25464 32419
rect 25412 32376 25464 32385
rect 26976 32419 27028 32428
rect 26976 32385 26985 32419
rect 26985 32385 27019 32419
rect 27019 32385 27028 32419
rect 26976 32376 27028 32385
rect 27068 32376 27120 32428
rect 12992 32240 13044 32292
rect 848 32172 900 32224
rect 11980 32215 12032 32224
rect 11980 32181 11989 32215
rect 11989 32181 12023 32215
rect 12023 32181 12032 32215
rect 11980 32172 12032 32181
rect 12440 32172 12492 32224
rect 13820 32172 13872 32224
rect 14004 32172 14056 32224
rect 17868 32172 17920 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 12992 32011 13044 32020
rect 12992 31977 13001 32011
rect 13001 31977 13035 32011
rect 13035 31977 13044 32011
rect 12992 31968 13044 31977
rect 13084 31968 13136 32020
rect 24400 32011 24452 32020
rect 24400 31977 24409 32011
rect 24409 31977 24443 32011
rect 24443 31977 24452 32011
rect 24400 31968 24452 31977
rect 24768 32011 24820 32020
rect 24768 31977 24777 32011
rect 24777 31977 24811 32011
rect 24811 31977 24820 32011
rect 24768 31968 24820 31977
rect 26148 31968 26200 32020
rect 27068 31968 27120 32020
rect 14188 31900 14240 31952
rect 848 31764 900 31816
rect 8852 31764 8904 31816
rect 11704 31807 11756 31816
rect 11704 31773 11713 31807
rect 11713 31773 11747 31807
rect 11747 31773 11756 31807
rect 11704 31764 11756 31773
rect 12716 31832 12768 31884
rect 12900 31764 12952 31816
rect 8668 31696 8720 31748
rect 10324 31671 10376 31680
rect 10324 31637 10333 31671
rect 10333 31637 10367 31671
rect 10367 31637 10376 31671
rect 10324 31628 10376 31637
rect 13360 31875 13412 31884
rect 13360 31841 13369 31875
rect 13369 31841 13403 31875
rect 13403 31841 13412 31875
rect 13360 31832 13412 31841
rect 14004 31832 14056 31884
rect 20904 31900 20956 31952
rect 21272 31900 21324 31952
rect 16304 31764 16356 31816
rect 16580 31764 16632 31816
rect 24308 31900 24360 31952
rect 24860 31900 24912 31952
rect 28448 31943 28500 31952
rect 28448 31909 28457 31943
rect 28457 31909 28491 31943
rect 28491 31909 28500 31943
rect 28448 31900 28500 31909
rect 24216 31807 24268 31816
rect 24216 31773 24225 31807
rect 24225 31773 24259 31807
rect 24259 31773 24268 31807
rect 24216 31764 24268 31773
rect 13544 31739 13596 31748
rect 13544 31705 13553 31739
rect 13553 31705 13587 31739
rect 13587 31705 13596 31739
rect 13544 31696 13596 31705
rect 13820 31696 13872 31748
rect 26056 31832 26108 31884
rect 26516 31875 26568 31884
rect 26516 31841 26525 31875
rect 26525 31841 26559 31875
rect 26559 31841 26568 31875
rect 26516 31832 26568 31841
rect 25688 31764 25740 31816
rect 26792 31807 26844 31816
rect 26792 31773 26801 31807
rect 26801 31773 26835 31807
rect 26835 31773 26844 31807
rect 26792 31764 26844 31773
rect 28356 31764 28408 31816
rect 25044 31696 25096 31748
rect 13268 31628 13320 31680
rect 24952 31628 25004 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 8668 31467 8720 31476
rect 8668 31433 8677 31467
rect 8677 31433 8711 31467
rect 8711 31433 8720 31467
rect 8668 31424 8720 31433
rect 12808 31424 12860 31476
rect 25412 31467 25464 31476
rect 25412 31433 25421 31467
rect 25421 31433 25455 31467
rect 25455 31433 25464 31467
rect 25412 31424 25464 31433
rect 6920 31288 6972 31340
rect 8576 31356 8628 31408
rect 11704 31288 11756 31340
rect 5816 31263 5868 31272
rect 5816 31229 5825 31263
rect 5825 31229 5859 31263
rect 5859 31229 5868 31263
rect 5816 31220 5868 31229
rect 6460 31220 6512 31272
rect 9220 31220 9272 31272
rect 11888 31331 11940 31340
rect 11888 31297 11897 31331
rect 11897 31297 11931 31331
rect 11931 31297 11940 31331
rect 11888 31288 11940 31297
rect 11980 31331 12032 31340
rect 11980 31297 11989 31331
rect 11989 31297 12023 31331
rect 12023 31297 12032 31331
rect 11980 31288 12032 31297
rect 12716 31356 12768 31408
rect 13084 31356 13136 31408
rect 12440 31288 12492 31340
rect 12624 31288 12676 31340
rect 12900 31288 12952 31340
rect 13176 31331 13228 31340
rect 13176 31297 13185 31331
rect 13185 31297 13219 31331
rect 13219 31297 13228 31331
rect 13176 31288 13228 31297
rect 24952 31331 25004 31340
rect 24952 31297 24961 31331
rect 24961 31297 24995 31331
rect 24995 31297 25004 31331
rect 24952 31288 25004 31297
rect 25044 31331 25096 31340
rect 25044 31297 25053 31331
rect 25053 31297 25087 31331
rect 25087 31297 25096 31331
rect 25044 31288 25096 31297
rect 25688 31331 25740 31340
rect 25688 31297 25697 31331
rect 25697 31297 25731 31331
rect 25731 31297 25740 31331
rect 25688 31288 25740 31297
rect 12624 31152 12676 31204
rect 12808 31152 12860 31204
rect 26148 31220 26200 31272
rect 5448 31127 5500 31136
rect 5448 31093 5457 31127
rect 5457 31093 5491 31127
rect 5491 31093 5500 31127
rect 5448 31084 5500 31093
rect 6368 31127 6420 31136
rect 6368 31093 6377 31127
rect 6377 31093 6411 31127
rect 6411 31093 6420 31127
rect 6368 31084 6420 31093
rect 11520 31127 11572 31136
rect 11520 31093 11529 31127
rect 11529 31093 11563 31127
rect 11563 31093 11572 31127
rect 11520 31084 11572 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 6460 30923 6512 30932
rect 6460 30889 6469 30923
rect 6469 30889 6503 30923
rect 6503 30889 6512 30923
rect 6460 30880 6512 30889
rect 12532 30880 12584 30932
rect 848 30744 900 30796
rect 2964 30676 3016 30728
rect 6920 30744 6972 30796
rect 7104 30787 7156 30796
rect 7104 30753 7113 30787
rect 7113 30753 7147 30787
rect 7147 30753 7156 30787
rect 7104 30744 7156 30753
rect 15660 30787 15712 30796
rect 15660 30753 15669 30787
rect 15669 30753 15703 30787
rect 15703 30753 15712 30787
rect 15660 30744 15712 30753
rect 6736 30676 6788 30728
rect 9588 30676 9640 30728
rect 11520 30719 11572 30728
rect 11520 30685 11554 30719
rect 11554 30685 11572 30719
rect 11520 30676 11572 30685
rect 12716 30719 12768 30728
rect 12716 30685 12725 30719
rect 12725 30685 12759 30719
rect 12759 30685 12768 30719
rect 12716 30676 12768 30685
rect 12900 30719 12952 30728
rect 12900 30685 12909 30719
rect 12909 30685 12943 30719
rect 12943 30685 12952 30719
rect 12900 30676 12952 30685
rect 15568 30719 15620 30728
rect 15568 30685 15577 30719
rect 15577 30685 15611 30719
rect 15611 30685 15620 30719
rect 15568 30676 15620 30685
rect 9220 30608 9272 30660
rect 6644 30540 6696 30592
rect 6920 30540 6972 30592
rect 8944 30540 8996 30592
rect 12624 30583 12676 30592
rect 12624 30549 12633 30583
rect 12633 30549 12667 30583
rect 12667 30549 12676 30583
rect 12624 30540 12676 30549
rect 13820 30540 13872 30592
rect 15108 30540 15160 30592
rect 15936 30583 15988 30592
rect 15936 30549 15945 30583
rect 15945 30549 15979 30583
rect 15979 30549 15988 30583
rect 15936 30540 15988 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 11888 30336 11940 30388
rect 13636 30336 13688 30388
rect 6644 30311 6696 30320
rect 4712 30132 4764 30184
rect 5448 30200 5500 30252
rect 6644 30277 6678 30311
rect 6678 30277 6696 30311
rect 6644 30268 6696 30277
rect 8852 30268 8904 30320
rect 9588 30268 9640 30320
rect 7012 30200 7064 30252
rect 7380 30200 7432 30252
rect 15936 30268 15988 30320
rect 7748 30107 7800 30116
rect 7748 30073 7757 30107
rect 7757 30073 7791 30107
rect 7791 30073 7800 30107
rect 7748 30064 7800 30073
rect 7104 29996 7156 30048
rect 7288 29996 7340 30048
rect 9220 29996 9272 30048
rect 15292 30243 15344 30252
rect 15292 30209 15301 30243
rect 15301 30209 15335 30243
rect 15335 30209 15344 30243
rect 15292 30200 15344 30209
rect 16304 30243 16356 30252
rect 16304 30209 16313 30243
rect 16313 30209 16347 30243
rect 16347 30209 16356 30243
rect 16304 30200 16356 30209
rect 16396 30200 16448 30252
rect 26976 30243 27028 30252
rect 26976 30209 26985 30243
rect 26985 30209 27019 30243
rect 27019 30209 27028 30243
rect 26976 30200 27028 30209
rect 27068 30200 27120 30252
rect 10692 30175 10744 30184
rect 10692 30141 10701 30175
rect 10701 30141 10735 30175
rect 10735 30141 10744 30175
rect 10692 30132 10744 30141
rect 12624 30132 12676 30184
rect 13544 30132 13596 30184
rect 15660 30175 15712 30184
rect 15660 30141 15669 30175
rect 15669 30141 15703 30175
rect 15703 30141 15712 30175
rect 15660 30132 15712 30141
rect 19340 30132 19392 30184
rect 28356 30107 28408 30116
rect 28356 30073 28365 30107
rect 28365 30073 28399 30107
rect 28399 30073 28408 30107
rect 28356 30064 28408 30073
rect 11336 29996 11388 30048
rect 16212 30039 16264 30048
rect 16212 30005 16221 30039
rect 16221 30005 16255 30039
rect 16255 30005 16264 30039
rect 16212 29996 16264 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 6828 29835 6880 29844
rect 6828 29801 6837 29835
rect 6837 29801 6871 29835
rect 6871 29801 6880 29835
rect 6828 29792 6880 29801
rect 6736 29767 6788 29776
rect 6736 29733 6745 29767
rect 6745 29733 6779 29767
rect 6779 29733 6788 29767
rect 6736 29724 6788 29733
rect 7748 29792 7800 29844
rect 11336 29835 11388 29844
rect 11336 29801 11345 29835
rect 11345 29801 11379 29835
rect 11379 29801 11388 29835
rect 11336 29792 11388 29801
rect 848 29588 900 29640
rect 2964 29631 3016 29640
rect 2964 29597 2973 29631
rect 2973 29597 3007 29631
rect 3007 29597 3016 29631
rect 2964 29588 3016 29597
rect 4712 29588 4764 29640
rect 7104 29631 7156 29640
rect 7104 29597 7113 29631
rect 7113 29597 7147 29631
rect 7147 29597 7156 29631
rect 7104 29588 7156 29597
rect 8944 29699 8996 29708
rect 8944 29665 8953 29699
rect 8953 29665 8987 29699
rect 8987 29665 8996 29699
rect 8944 29656 8996 29665
rect 10600 29656 10652 29708
rect 17776 29656 17828 29708
rect 8852 29588 8904 29640
rect 9496 29588 9548 29640
rect 10416 29631 10468 29640
rect 10416 29597 10425 29631
rect 10425 29597 10459 29631
rect 10459 29597 10468 29631
rect 10416 29588 10468 29597
rect 12348 29588 12400 29640
rect 16212 29588 16264 29640
rect 6368 29520 6420 29572
rect 6736 29520 6788 29572
rect 7656 29563 7708 29572
rect 7656 29529 7679 29563
rect 7679 29529 7708 29563
rect 7656 29520 7708 29529
rect 8668 29452 8720 29504
rect 10324 29520 10376 29572
rect 9404 29452 9456 29504
rect 9680 29495 9732 29504
rect 9680 29461 9689 29495
rect 9689 29461 9723 29495
rect 9723 29461 9732 29495
rect 9680 29452 9732 29461
rect 10692 29452 10744 29504
rect 15292 29452 15344 29504
rect 16304 29452 16356 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 5816 29248 5868 29300
rect 7656 29248 7708 29300
rect 9680 29248 9732 29300
rect 10416 29248 10468 29300
rect 6920 29112 6972 29164
rect 7288 29155 7340 29164
rect 7288 29121 7297 29155
rect 7297 29121 7331 29155
rect 7331 29121 7340 29155
rect 7288 29112 7340 29121
rect 7380 29155 7432 29164
rect 7380 29121 7389 29155
rect 7389 29121 7423 29155
rect 7423 29121 7432 29155
rect 7380 29112 7432 29121
rect 9220 29180 9272 29232
rect 8576 29155 8628 29164
rect 8576 29121 8585 29155
rect 8585 29121 8619 29155
rect 8619 29121 8628 29155
rect 8576 29112 8628 29121
rect 8852 29155 8904 29164
rect 8852 29121 8861 29155
rect 8861 29121 8895 29155
rect 8895 29121 8904 29155
rect 8852 29112 8904 29121
rect 8668 29044 8720 29096
rect 10600 29155 10652 29164
rect 10600 29121 10609 29155
rect 10609 29121 10643 29155
rect 10643 29121 10652 29155
rect 10600 29112 10652 29121
rect 15108 29155 15160 29164
rect 15108 29121 15117 29155
rect 15117 29121 15151 29155
rect 15151 29121 15160 29155
rect 15108 29112 15160 29121
rect 18328 29155 18380 29164
rect 18328 29121 18337 29155
rect 18337 29121 18371 29155
rect 18371 29121 18380 29155
rect 18328 29112 18380 29121
rect 18420 29155 18472 29164
rect 18420 29121 18429 29155
rect 18429 29121 18463 29155
rect 18463 29121 18472 29155
rect 18420 29112 18472 29121
rect 19340 29112 19392 29164
rect 19984 29112 20036 29164
rect 848 28976 900 29028
rect 17500 28976 17552 29028
rect 27068 28976 27120 29028
rect 10324 28951 10376 28960
rect 10324 28917 10333 28951
rect 10333 28917 10367 28951
rect 10367 28917 10376 28951
rect 10324 28908 10376 28917
rect 10784 28951 10836 28960
rect 10784 28917 10793 28951
rect 10793 28917 10827 28951
rect 10827 28917 10836 28951
rect 10784 28908 10836 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 18420 28747 18472 28756
rect 18420 28713 18429 28747
rect 18429 28713 18463 28747
rect 18463 28713 18472 28747
rect 18420 28704 18472 28713
rect 22376 28636 22428 28688
rect 17592 28568 17644 28620
rect 9404 28500 9456 28552
rect 9496 28543 9548 28552
rect 9496 28509 9505 28543
rect 9505 28509 9539 28543
rect 9539 28509 9548 28543
rect 9496 28500 9548 28509
rect 8944 28407 8996 28416
rect 8944 28373 8953 28407
rect 8953 28373 8987 28407
rect 8987 28373 8996 28407
rect 8944 28364 8996 28373
rect 10784 28432 10836 28484
rect 16304 28432 16356 28484
rect 17868 28543 17920 28552
rect 17868 28509 17877 28543
rect 17877 28509 17911 28543
rect 17911 28509 17920 28543
rect 17868 28500 17920 28509
rect 19432 28568 19484 28620
rect 18236 28543 18288 28552
rect 18236 28509 18245 28543
rect 18245 28509 18279 28543
rect 18279 28509 18288 28543
rect 18236 28500 18288 28509
rect 10692 28364 10744 28416
rect 17592 28407 17644 28416
rect 17592 28373 17601 28407
rect 17601 28373 17635 28407
rect 17635 28373 17644 28407
rect 17592 28364 17644 28373
rect 17960 28432 18012 28484
rect 19800 28543 19852 28552
rect 19800 28509 19809 28543
rect 19809 28509 19843 28543
rect 19843 28509 19852 28543
rect 19800 28500 19852 28509
rect 19984 28543 20036 28552
rect 19984 28509 19993 28543
rect 19993 28509 20027 28543
rect 20027 28509 20036 28543
rect 19984 28500 20036 28509
rect 20904 28543 20956 28552
rect 20904 28509 20913 28543
rect 20913 28509 20947 28543
rect 20947 28509 20956 28543
rect 20904 28500 20956 28509
rect 20260 28432 20312 28484
rect 21272 28500 21324 28552
rect 19340 28364 19392 28416
rect 20812 28364 20864 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 18328 28160 18380 28212
rect 19432 28203 19484 28212
rect 19432 28169 19441 28203
rect 19441 28169 19475 28203
rect 19475 28169 19484 28203
rect 19432 28160 19484 28169
rect 17684 28092 17736 28144
rect 17132 28024 17184 28076
rect 17592 28067 17644 28076
rect 17592 28033 17602 28067
rect 17602 28033 17636 28067
rect 17636 28033 17644 28067
rect 17592 28024 17644 28033
rect 22008 28092 22060 28144
rect 19616 28024 19668 28076
rect 18144 27956 18196 28008
rect 21180 28024 21232 28076
rect 28540 27931 28592 27940
rect 28540 27897 28549 27931
rect 28549 27897 28583 27931
rect 28583 27897 28592 27931
rect 28540 27888 28592 27897
rect 21548 27863 21600 27872
rect 21548 27829 21557 27863
rect 21557 27829 21591 27863
rect 21591 27829 21600 27863
rect 21548 27820 21600 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 16764 27548 16816 27600
rect 18236 27616 18288 27668
rect 19708 27616 19760 27668
rect 18144 27591 18196 27600
rect 18144 27557 18153 27591
rect 18153 27557 18187 27591
rect 18187 27557 18196 27591
rect 18144 27548 18196 27557
rect 19340 27548 19392 27600
rect 20904 27616 20956 27668
rect 13452 27455 13504 27464
rect 13452 27421 13461 27455
rect 13461 27421 13495 27455
rect 13495 27421 13504 27455
rect 13452 27412 13504 27421
rect 13636 27455 13688 27464
rect 13636 27421 13645 27455
rect 13645 27421 13679 27455
rect 13679 27421 13688 27455
rect 13636 27412 13688 27421
rect 17592 27455 17644 27464
rect 17592 27421 17601 27455
rect 17601 27421 17635 27455
rect 17635 27421 17644 27455
rect 17592 27412 17644 27421
rect 17868 27455 17920 27464
rect 17868 27421 17877 27455
rect 17877 27421 17911 27455
rect 17911 27421 17920 27455
rect 17868 27412 17920 27421
rect 17960 27455 18012 27464
rect 17960 27421 17969 27455
rect 17969 27421 18003 27455
rect 18003 27421 18012 27455
rect 17960 27412 18012 27421
rect 18972 27455 19024 27464
rect 18972 27421 18981 27455
rect 18981 27421 19015 27455
rect 19015 27421 19024 27455
rect 18972 27412 19024 27421
rect 19064 27455 19116 27464
rect 19064 27421 19073 27455
rect 19073 27421 19107 27455
rect 19107 27421 19116 27455
rect 19064 27412 19116 27421
rect 16304 27344 16356 27396
rect 17684 27344 17736 27396
rect 20812 27455 20864 27464
rect 20812 27421 20821 27455
rect 20821 27421 20855 27455
rect 20855 27421 20864 27455
rect 20812 27412 20864 27421
rect 21548 27523 21600 27532
rect 21548 27489 21557 27523
rect 21557 27489 21591 27523
rect 21591 27489 21600 27523
rect 21548 27480 21600 27489
rect 22008 27523 22060 27532
rect 22008 27489 22017 27523
rect 22017 27489 22051 27523
rect 22051 27489 22060 27523
rect 22008 27480 22060 27489
rect 21824 27455 21876 27464
rect 21824 27421 21833 27455
rect 21833 27421 21867 27455
rect 21867 27421 21876 27455
rect 21824 27412 21876 27421
rect 22376 27455 22428 27464
rect 22376 27421 22385 27455
rect 22385 27421 22419 27455
rect 22419 27421 22428 27455
rect 22376 27412 22428 27421
rect 21180 27344 21232 27396
rect 21548 27344 21600 27396
rect 14004 27276 14056 27328
rect 17132 27319 17184 27328
rect 17132 27285 17141 27319
rect 17141 27285 17175 27319
rect 17175 27285 17184 27319
rect 17132 27276 17184 27285
rect 19984 27276 20036 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 12900 27072 12952 27124
rect 17684 27115 17736 27124
rect 17684 27081 17693 27115
rect 17693 27081 17727 27115
rect 17727 27081 17736 27115
rect 17684 27072 17736 27081
rect 19064 27115 19116 27124
rect 19064 27081 19073 27115
rect 19073 27081 19107 27115
rect 19107 27081 19116 27115
rect 19064 27072 19116 27081
rect 8944 27004 8996 27056
rect 16948 27004 17000 27056
rect 17500 27047 17552 27056
rect 17500 27013 17509 27047
rect 17509 27013 17543 27047
rect 17543 27013 17552 27047
rect 17500 27004 17552 27013
rect 21548 27004 21600 27056
rect 12992 26936 13044 26988
rect 13820 26979 13872 26988
rect 13820 26945 13829 26979
rect 13829 26945 13863 26979
rect 13863 26945 13872 26979
rect 13820 26936 13872 26945
rect 14004 26979 14056 26988
rect 14004 26945 14013 26979
rect 14013 26945 14047 26979
rect 14047 26945 14056 26979
rect 14004 26936 14056 26945
rect 8944 26911 8996 26920
rect 8944 26877 8953 26911
rect 8953 26877 8987 26911
rect 8987 26877 8996 26911
rect 8944 26868 8996 26877
rect 12624 26911 12676 26920
rect 12624 26877 12633 26911
rect 12633 26877 12667 26911
rect 12667 26877 12676 26911
rect 12624 26868 12676 26877
rect 13176 26800 13228 26852
rect 13636 26911 13688 26920
rect 13636 26877 13645 26911
rect 13645 26877 13679 26911
rect 13679 26877 13688 26911
rect 13636 26868 13688 26877
rect 13728 26868 13780 26920
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 16856 26936 16908 26988
rect 17960 26936 18012 26988
rect 19248 26936 19300 26988
rect 19984 26936 20036 26988
rect 21180 26979 21232 26988
rect 21180 26945 21189 26979
rect 21189 26945 21223 26979
rect 21223 26945 21232 26979
rect 21180 26936 21232 26945
rect 18236 26800 18288 26852
rect 10324 26775 10376 26784
rect 10324 26741 10333 26775
rect 10333 26741 10367 26775
rect 10367 26741 10376 26775
rect 10324 26732 10376 26741
rect 13084 26775 13136 26784
rect 13084 26741 13093 26775
rect 13093 26741 13127 26775
rect 13127 26741 13136 26775
rect 13084 26732 13136 26741
rect 14464 26775 14516 26784
rect 14464 26741 14473 26775
rect 14473 26741 14507 26775
rect 14507 26741 14516 26775
rect 14464 26732 14516 26741
rect 20812 26732 20864 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 13636 26528 13688 26580
rect 14188 26528 14240 26580
rect 13912 26460 13964 26512
rect 16672 26571 16724 26580
rect 16672 26537 16681 26571
rect 16681 26537 16715 26571
rect 16715 26537 16724 26571
rect 16672 26528 16724 26537
rect 19892 26528 19944 26580
rect 19984 26571 20036 26580
rect 19984 26537 19993 26571
rect 19993 26537 20027 26571
rect 20027 26537 20036 26571
rect 19984 26528 20036 26537
rect 21824 26528 21876 26580
rect 17868 26460 17920 26512
rect 19800 26460 19852 26512
rect 8944 26392 8996 26444
rect 12624 26324 12676 26376
rect 14188 26324 14240 26376
rect 14372 26367 14424 26376
rect 14372 26333 14381 26367
rect 14381 26333 14415 26367
rect 14415 26333 14424 26367
rect 14372 26324 14424 26333
rect 14464 26324 14516 26376
rect 24492 26392 24544 26444
rect 19248 26324 19300 26376
rect 12256 26299 12308 26308
rect 12256 26265 12290 26299
rect 12290 26265 12308 26299
rect 12256 26256 12308 26265
rect 18972 26256 19024 26308
rect 19616 26256 19668 26308
rect 20260 26367 20312 26376
rect 20260 26333 20269 26367
rect 20269 26333 20303 26367
rect 20303 26333 20312 26367
rect 20260 26324 20312 26333
rect 20904 26324 20956 26376
rect 12348 26188 12400 26240
rect 12992 26188 13044 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 9496 25984 9548 26036
rect 12256 26027 12308 26036
rect 12256 25993 12265 26027
rect 12265 25993 12299 26027
rect 12299 25993 12308 26027
rect 12256 25984 12308 25993
rect 13176 25984 13228 26036
rect 13452 25984 13504 26036
rect 17592 25984 17644 26036
rect 9404 25891 9456 25900
rect 9404 25857 9413 25891
rect 9413 25857 9447 25891
rect 9447 25857 9456 25891
rect 9404 25848 9456 25857
rect 9864 25848 9916 25900
rect 10324 25848 10376 25900
rect 12440 25848 12492 25900
rect 12256 25780 12308 25832
rect 12348 25780 12400 25832
rect 12624 25891 12676 25900
rect 12624 25857 12633 25891
rect 12633 25857 12667 25891
rect 12667 25857 12676 25891
rect 12624 25848 12676 25857
rect 12900 25891 12952 25900
rect 12900 25857 12909 25891
rect 12909 25857 12943 25891
rect 12943 25857 12952 25891
rect 12900 25848 12952 25857
rect 12992 25848 13044 25900
rect 13084 25823 13136 25832
rect 13084 25789 13093 25823
rect 13093 25789 13127 25823
rect 13127 25789 13136 25823
rect 13084 25780 13136 25789
rect 16120 25891 16172 25900
rect 16120 25857 16129 25891
rect 16129 25857 16163 25891
rect 16163 25857 16172 25891
rect 16120 25848 16172 25857
rect 16764 25916 16816 25968
rect 16948 25959 17000 25968
rect 16948 25925 16957 25959
rect 16957 25925 16991 25959
rect 16991 25925 17000 25959
rect 16948 25916 17000 25925
rect 16304 25891 16356 25900
rect 16304 25857 16313 25891
rect 16313 25857 16347 25891
rect 16347 25857 16356 25891
rect 16304 25848 16356 25857
rect 16856 25891 16908 25900
rect 16856 25857 16860 25891
rect 16860 25857 16894 25891
rect 16894 25857 16908 25891
rect 16856 25848 16908 25857
rect 17224 25891 17276 25900
rect 17224 25857 17232 25891
rect 17232 25857 17266 25891
rect 17266 25857 17276 25891
rect 17224 25848 17276 25857
rect 13728 25780 13780 25832
rect 17868 25891 17920 25900
rect 17868 25857 17877 25891
rect 17877 25857 17911 25891
rect 17911 25857 17920 25891
rect 17868 25848 17920 25857
rect 19432 25712 19484 25764
rect 12164 25687 12216 25696
rect 12164 25653 12173 25687
rect 12173 25653 12207 25687
rect 12207 25653 12216 25687
rect 12164 25644 12216 25653
rect 12624 25644 12676 25696
rect 13636 25644 13688 25696
rect 13728 25687 13780 25696
rect 13728 25653 13737 25687
rect 13737 25653 13771 25687
rect 13771 25653 13780 25687
rect 13728 25644 13780 25653
rect 15936 25687 15988 25696
rect 15936 25653 15945 25687
rect 15945 25653 15979 25687
rect 15979 25653 15988 25687
rect 15936 25644 15988 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 13728 25440 13780 25492
rect 12992 25415 13044 25424
rect 12992 25381 13001 25415
rect 13001 25381 13035 25415
rect 13035 25381 13044 25415
rect 12992 25372 13044 25381
rect 13176 25372 13228 25424
rect 13636 25372 13688 25424
rect 8392 25304 8444 25356
rect 8760 25304 8812 25356
rect 12164 25304 12216 25356
rect 7012 25279 7064 25288
rect 7012 25245 7021 25279
rect 7021 25245 7055 25279
rect 7055 25245 7064 25279
rect 7012 25236 7064 25245
rect 12256 25279 12308 25288
rect 12256 25245 12265 25279
rect 12265 25245 12299 25279
rect 12299 25245 12308 25279
rect 12256 25236 12308 25245
rect 12440 25279 12492 25288
rect 12440 25245 12449 25279
rect 12449 25245 12483 25279
rect 12483 25245 12492 25279
rect 12440 25236 12492 25245
rect 12532 25279 12584 25288
rect 12532 25245 12541 25279
rect 12541 25245 12575 25279
rect 12575 25245 12584 25279
rect 12532 25236 12584 25245
rect 12900 25304 12952 25356
rect 13820 25304 13872 25356
rect 13268 25236 13320 25288
rect 15384 25236 15436 25288
rect 16120 25236 16172 25288
rect 17132 25236 17184 25288
rect 7840 25168 7892 25220
rect 6368 25100 6420 25152
rect 8116 25100 8168 25152
rect 12348 25100 12400 25152
rect 13912 25168 13964 25220
rect 15660 25100 15712 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 12532 24896 12584 24948
rect 13544 24896 13596 24948
rect 848 24760 900 24812
rect 2504 24735 2556 24744
rect 2504 24701 2513 24735
rect 2513 24701 2547 24735
rect 2547 24701 2556 24735
rect 2504 24692 2556 24701
rect 9496 24828 9548 24880
rect 16856 24828 16908 24880
rect 19616 24828 19668 24880
rect 4712 24803 4764 24812
rect 4712 24769 4721 24803
rect 4721 24769 4755 24803
rect 4755 24769 4764 24803
rect 4712 24760 4764 24769
rect 4804 24760 4856 24812
rect 7472 24803 7524 24812
rect 7472 24769 7490 24803
rect 7490 24769 7524 24803
rect 7472 24760 7524 24769
rect 13360 24760 13412 24812
rect 13912 24803 13964 24812
rect 13912 24769 13921 24803
rect 13921 24769 13955 24803
rect 13955 24769 13964 24803
rect 13912 24760 13964 24769
rect 8392 24692 8444 24744
rect 13636 24624 13688 24676
rect 5448 24556 5500 24608
rect 6092 24599 6144 24608
rect 6092 24565 6101 24599
rect 6101 24565 6135 24599
rect 6135 24565 6144 24599
rect 6092 24556 6144 24565
rect 7012 24556 7064 24608
rect 10140 24599 10192 24608
rect 10140 24565 10149 24599
rect 10149 24565 10183 24599
rect 10183 24565 10192 24599
rect 10140 24556 10192 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 4804 24395 4856 24404
rect 4804 24361 4813 24395
rect 4813 24361 4847 24395
rect 4847 24361 4856 24395
rect 4804 24352 4856 24361
rect 5448 24352 5500 24404
rect 6736 24352 6788 24404
rect 7840 24395 7892 24404
rect 7840 24361 7849 24395
rect 7849 24361 7883 24395
rect 7883 24361 7892 24395
rect 7840 24352 7892 24361
rect 6368 24284 6420 24336
rect 5448 24259 5500 24268
rect 5448 24225 5457 24259
rect 5457 24225 5491 24259
rect 5491 24225 5500 24259
rect 5448 24216 5500 24225
rect 6092 24216 6144 24268
rect 12440 24284 12492 24336
rect 2504 24148 2556 24200
rect 5908 24148 5960 24200
rect 6368 24191 6420 24200
rect 6368 24157 6377 24191
rect 6377 24157 6411 24191
rect 6411 24157 6420 24191
rect 6368 24148 6420 24157
rect 8300 24216 8352 24268
rect 9404 24216 9456 24268
rect 13544 24259 13596 24268
rect 13544 24225 13553 24259
rect 13553 24225 13587 24259
rect 13587 24225 13596 24259
rect 13544 24216 13596 24225
rect 8116 24191 8168 24200
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 13636 24191 13688 24200
rect 13636 24157 13645 24191
rect 13645 24157 13679 24191
rect 13679 24157 13688 24191
rect 13636 24148 13688 24157
rect 7012 24080 7064 24132
rect 7288 24123 7340 24132
rect 7288 24089 7297 24123
rect 7297 24089 7331 24123
rect 7331 24089 7340 24123
rect 7288 24080 7340 24089
rect 6000 24012 6052 24064
rect 7196 24055 7248 24064
rect 7196 24021 7205 24055
rect 7205 24021 7239 24055
rect 7239 24021 7248 24055
rect 7196 24012 7248 24021
rect 7748 24055 7800 24064
rect 7748 24021 7757 24055
rect 7757 24021 7791 24055
rect 7791 24021 7800 24055
rect 7748 24012 7800 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 6368 23808 6420 23860
rect 7472 23851 7524 23860
rect 7472 23817 7481 23851
rect 7481 23817 7515 23851
rect 7515 23817 7524 23851
rect 7472 23808 7524 23817
rect 10140 23740 10192 23792
rect 5908 23715 5960 23724
rect 5908 23681 5917 23715
rect 5917 23681 5951 23715
rect 5951 23681 5960 23715
rect 5908 23672 5960 23681
rect 6000 23715 6052 23724
rect 6000 23681 6009 23715
rect 6009 23681 6043 23715
rect 6043 23681 6052 23715
rect 6000 23672 6052 23681
rect 6736 23715 6788 23724
rect 6736 23681 6745 23715
rect 6745 23681 6779 23715
rect 6779 23681 6788 23715
rect 6736 23672 6788 23681
rect 7196 23715 7248 23724
rect 7196 23681 7205 23715
rect 7205 23681 7239 23715
rect 7239 23681 7248 23715
rect 7196 23672 7248 23681
rect 6368 23647 6420 23656
rect 6368 23613 6377 23647
rect 6377 23613 6411 23647
rect 6411 23613 6420 23647
rect 6368 23604 6420 23613
rect 6828 23647 6880 23656
rect 6828 23613 6837 23647
rect 6837 23613 6871 23647
rect 6871 23613 6880 23647
rect 6828 23604 6880 23613
rect 8300 23672 8352 23724
rect 9772 23715 9824 23724
rect 9772 23681 9781 23715
rect 9781 23681 9815 23715
rect 9815 23681 9824 23715
rect 9772 23672 9824 23681
rect 10416 23715 10468 23724
rect 10416 23681 10425 23715
rect 10425 23681 10459 23715
rect 10459 23681 10468 23715
rect 10416 23672 10468 23681
rect 13636 23672 13688 23724
rect 9864 23647 9916 23656
rect 9864 23613 9873 23647
rect 9873 23613 9907 23647
rect 9907 23613 9916 23647
rect 9864 23604 9916 23613
rect 11428 23536 11480 23588
rect 15292 23715 15344 23724
rect 15292 23681 15301 23715
rect 15301 23681 15335 23715
rect 15335 23681 15344 23715
rect 15292 23672 15344 23681
rect 15660 23715 15712 23724
rect 15660 23681 15669 23715
rect 15669 23681 15703 23715
rect 15703 23681 15712 23715
rect 15660 23672 15712 23681
rect 15752 23715 15804 23724
rect 15752 23681 15762 23715
rect 15762 23681 15796 23715
rect 15796 23681 15804 23715
rect 15752 23672 15804 23681
rect 15936 23783 15988 23792
rect 15936 23749 15945 23783
rect 15945 23749 15979 23783
rect 15979 23749 15988 23783
rect 15936 23740 15988 23749
rect 17224 23851 17276 23860
rect 17224 23817 17233 23851
rect 17233 23817 17267 23851
rect 17267 23817 17276 23851
rect 17224 23808 17276 23817
rect 18972 23808 19024 23860
rect 18144 23740 18196 23792
rect 19616 23783 19668 23792
rect 19616 23749 19625 23783
rect 19625 23749 19659 23783
rect 19659 23749 19668 23783
rect 19616 23740 19668 23749
rect 16120 23715 16172 23724
rect 16120 23681 16134 23715
rect 16134 23681 16168 23715
rect 16168 23681 16172 23715
rect 16120 23672 16172 23681
rect 5724 23511 5776 23520
rect 5724 23477 5733 23511
rect 5733 23477 5767 23511
rect 5767 23477 5776 23511
rect 5724 23468 5776 23477
rect 7104 23468 7156 23520
rect 11244 23468 11296 23520
rect 16856 23468 16908 23520
rect 17960 23604 18012 23656
rect 18972 23604 19024 23656
rect 28264 23715 28316 23724
rect 28264 23681 28273 23715
rect 28273 23681 28307 23715
rect 28307 23681 28316 23715
rect 28264 23672 28316 23681
rect 19432 23511 19484 23520
rect 19432 23477 19441 23511
rect 19441 23477 19475 23511
rect 19475 23477 19484 23511
rect 19432 23468 19484 23477
rect 19708 23511 19760 23520
rect 19708 23477 19717 23511
rect 19717 23477 19751 23511
rect 19751 23477 19760 23511
rect 19708 23468 19760 23477
rect 28448 23511 28500 23520
rect 28448 23477 28457 23511
rect 28457 23477 28491 23511
rect 28491 23477 28500 23511
rect 28448 23468 28500 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 10416 23264 10468 23316
rect 4712 23128 4764 23180
rect 5356 23060 5408 23112
rect 6828 23060 6880 23112
rect 7104 23103 7156 23112
rect 7104 23069 7113 23103
rect 7113 23069 7147 23103
rect 7147 23069 7156 23103
rect 7104 23060 7156 23069
rect 9956 23128 10008 23180
rect 13268 23264 13320 23316
rect 16856 23307 16908 23316
rect 16856 23273 16865 23307
rect 16865 23273 16899 23307
rect 16899 23273 16908 23307
rect 16856 23264 16908 23273
rect 28264 23264 28316 23316
rect 13360 23196 13412 23248
rect 8392 23060 8444 23112
rect 8944 23103 8996 23112
rect 8944 23069 8953 23103
rect 8953 23069 8987 23103
rect 8987 23069 8996 23103
rect 8944 23060 8996 23069
rect 9772 23060 9824 23112
rect 10600 23060 10652 23112
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 11428 23103 11480 23112
rect 11428 23069 11437 23103
rect 11437 23069 11471 23103
rect 11471 23069 11480 23103
rect 11428 23060 11480 23069
rect 18144 23196 18196 23248
rect 19616 23196 19668 23248
rect 17960 23128 18012 23180
rect 5724 22992 5776 23044
rect 6736 22924 6788 22976
rect 7012 23035 7064 23044
rect 7012 23001 7021 23035
rect 7021 23001 7055 23035
rect 7055 23001 7064 23035
rect 7012 22992 7064 23001
rect 8116 22992 8168 23044
rect 8668 22992 8720 23044
rect 10140 22992 10192 23044
rect 11704 23035 11756 23044
rect 11704 23001 11713 23035
rect 11713 23001 11747 23035
rect 11747 23001 11756 23035
rect 11704 22992 11756 23001
rect 7104 22924 7156 22976
rect 7472 22924 7524 22976
rect 8760 22967 8812 22976
rect 8760 22933 8769 22967
rect 8769 22933 8803 22967
rect 8803 22933 8812 22967
rect 8760 22924 8812 22933
rect 11796 22924 11848 22976
rect 15752 22992 15804 23044
rect 16764 22992 16816 23044
rect 18880 23103 18932 23112
rect 18880 23069 18889 23103
rect 18889 23069 18923 23103
rect 18923 23069 18932 23103
rect 18880 23060 18932 23069
rect 19432 23060 19484 23112
rect 27528 23103 27580 23112
rect 27528 23069 27537 23103
rect 27537 23069 27571 23103
rect 27571 23069 27580 23103
rect 27528 23060 27580 23069
rect 19708 22992 19760 23044
rect 12348 22967 12400 22976
rect 12348 22933 12357 22967
rect 12357 22933 12391 22967
rect 12391 22933 12400 22967
rect 12348 22924 12400 22933
rect 16120 22924 16172 22976
rect 17132 22967 17184 22976
rect 17132 22933 17141 22967
rect 17141 22933 17175 22967
rect 17175 22933 17184 22967
rect 17132 22924 17184 22933
rect 18512 22967 18564 22976
rect 18512 22933 18521 22967
rect 18521 22933 18555 22967
rect 18555 22933 18564 22967
rect 18512 22924 18564 22933
rect 19248 22967 19300 22976
rect 19248 22933 19257 22967
rect 19257 22933 19291 22967
rect 19291 22933 19300 22967
rect 19248 22924 19300 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 6368 22763 6420 22772
rect 6368 22729 6377 22763
rect 6377 22729 6411 22763
rect 6411 22729 6420 22763
rect 6368 22720 6420 22729
rect 6736 22763 6788 22772
rect 6736 22729 6745 22763
rect 6745 22729 6779 22763
rect 6779 22729 6788 22763
rect 6736 22720 6788 22729
rect 6920 22720 6972 22772
rect 8116 22763 8168 22772
rect 8116 22729 8125 22763
rect 8125 22729 8159 22763
rect 8159 22729 8168 22763
rect 8116 22720 8168 22729
rect 10600 22763 10652 22772
rect 10600 22729 10609 22763
rect 10609 22729 10643 22763
rect 10643 22729 10652 22763
rect 10600 22720 10652 22729
rect 15292 22720 15344 22772
rect 15752 22720 15804 22772
rect 16028 22720 16080 22772
rect 6828 22652 6880 22704
rect 8668 22695 8720 22704
rect 8668 22661 8677 22695
rect 8677 22661 8711 22695
rect 8711 22661 8720 22695
rect 8668 22652 8720 22661
rect 8760 22652 8812 22704
rect 6736 22584 6788 22636
rect 7288 22584 7340 22636
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 8300 22584 8352 22636
rect 9772 22584 9824 22636
rect 9956 22627 10008 22636
rect 9956 22593 9965 22627
rect 9965 22593 9999 22627
rect 9999 22593 10008 22627
rect 9956 22584 10008 22593
rect 10140 22627 10192 22636
rect 10140 22593 10149 22627
rect 10149 22593 10183 22627
rect 10183 22593 10192 22627
rect 10140 22584 10192 22593
rect 10508 22584 10560 22636
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 16120 22627 16172 22636
rect 16120 22593 16129 22627
rect 16129 22593 16163 22627
rect 16163 22593 16172 22627
rect 16120 22584 16172 22593
rect 16856 22584 16908 22636
rect 19248 22720 19300 22772
rect 19432 22720 19484 22772
rect 17960 22627 18012 22636
rect 17960 22593 17969 22627
rect 17969 22593 18003 22627
rect 18003 22593 18012 22627
rect 17960 22584 18012 22593
rect 18052 22584 18104 22636
rect 18512 22627 18564 22636
rect 18512 22593 18546 22627
rect 18546 22593 18564 22627
rect 18512 22584 18564 22593
rect 6828 22516 6880 22568
rect 11704 22516 11756 22568
rect 16580 22516 16632 22568
rect 18144 22516 18196 22568
rect 16764 22448 16816 22500
rect 28540 22559 28592 22568
rect 28540 22525 28549 22559
rect 28549 22525 28583 22559
rect 28583 22525 28592 22559
rect 28540 22516 28592 22525
rect 19616 22491 19668 22500
rect 19616 22457 19625 22491
rect 19625 22457 19659 22491
rect 19659 22457 19668 22491
rect 19616 22448 19668 22457
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 12348 22176 12400 22228
rect 6828 22108 6880 22160
rect 7104 22151 7156 22160
rect 7104 22117 7113 22151
rect 7113 22117 7147 22151
rect 7147 22117 7156 22151
rect 7104 22108 7156 22117
rect 18144 22176 18196 22228
rect 18604 22176 18656 22228
rect 18880 22176 18932 22228
rect 6920 22083 6972 22092
rect 6920 22049 6929 22083
rect 6929 22049 6963 22083
rect 6963 22049 6972 22083
rect 6920 22040 6972 22049
rect 11796 22040 11848 22092
rect 6736 21904 6788 21956
rect 7748 21972 7800 22024
rect 12440 22015 12492 22024
rect 6368 21879 6420 21888
rect 6368 21845 6377 21879
rect 6377 21845 6411 21879
rect 6411 21845 6420 21879
rect 6368 21836 6420 21845
rect 12440 21981 12449 22015
rect 12449 21981 12483 22015
rect 12483 21981 12492 22015
rect 12440 21972 12492 21981
rect 12532 21972 12584 22024
rect 19432 22040 19484 22092
rect 12256 21947 12308 21956
rect 12256 21913 12265 21947
rect 12265 21913 12299 21947
rect 12299 21913 12308 21947
rect 12256 21904 12308 21913
rect 12348 21904 12400 21956
rect 12992 21972 13044 22024
rect 17132 22015 17184 22024
rect 17132 21981 17150 22015
rect 17150 21981 17184 22015
rect 17132 21972 17184 21981
rect 17408 22015 17460 22024
rect 17408 21981 17417 22015
rect 17417 21981 17451 22015
rect 17451 21981 17460 22015
rect 17408 21972 17460 21981
rect 18052 21972 18104 22024
rect 18604 21972 18656 22024
rect 18788 22015 18840 22024
rect 18788 21981 18797 22015
rect 18797 21981 18831 22015
rect 18831 21981 18840 22015
rect 18788 21972 18840 21981
rect 18972 22015 19024 22024
rect 18972 21981 18981 22015
rect 18981 21981 19015 22015
rect 19015 21981 19024 22015
rect 18972 21972 19024 21981
rect 13820 21904 13872 21956
rect 14648 21904 14700 21956
rect 17960 21904 18012 21956
rect 12992 21836 13044 21888
rect 16580 21836 16632 21888
rect 18512 21836 18564 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 12440 21564 12492 21616
rect 12992 21360 13044 21412
rect 12164 21335 12216 21344
rect 12164 21301 12173 21335
rect 12173 21301 12207 21335
rect 12207 21301 12216 21335
rect 12164 21292 12216 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 7012 21088 7064 21140
rect 7196 21088 7248 21140
rect 7012 20927 7064 20936
rect 7012 20893 7021 20927
rect 7021 20893 7055 20927
rect 7055 20893 7064 20927
rect 7012 20884 7064 20893
rect 12440 20884 12492 20936
rect 12900 20884 12952 20936
rect 13176 20884 13228 20936
rect 8300 20816 8352 20868
rect 12992 20791 13044 20800
rect 12992 20757 13001 20791
rect 13001 20757 13035 20791
rect 13035 20757 13044 20791
rect 12992 20748 13044 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 16672 20544 16724 20596
rect 9496 20519 9548 20528
rect 9496 20485 9505 20519
rect 9505 20485 9539 20519
rect 9539 20485 9548 20519
rect 9496 20476 9548 20485
rect 6368 20408 6420 20460
rect 13820 20476 13872 20528
rect 14372 20476 14424 20528
rect 17408 20476 17460 20528
rect 7380 20340 7432 20392
rect 8208 20340 8260 20392
rect 12164 20383 12216 20392
rect 12164 20349 12173 20383
rect 12173 20349 12207 20383
rect 12207 20349 12216 20383
rect 12164 20340 12216 20349
rect 12900 20451 12952 20460
rect 12900 20417 12909 20451
rect 12909 20417 12943 20451
rect 12943 20417 12952 20451
rect 12900 20408 12952 20417
rect 12992 20451 13044 20460
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 12992 20408 13044 20417
rect 13084 20408 13136 20460
rect 13268 20408 13320 20460
rect 14464 20451 14516 20460
rect 14464 20417 14482 20451
rect 14482 20417 14516 20451
rect 14464 20408 14516 20417
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 14832 20451 14884 20460
rect 14832 20417 14841 20451
rect 14841 20417 14875 20451
rect 14875 20417 14884 20451
rect 14832 20408 14884 20417
rect 12532 20340 12584 20392
rect 15936 20408 15988 20460
rect 16028 20451 16080 20460
rect 16028 20417 16037 20451
rect 16037 20417 16071 20451
rect 16071 20417 16080 20451
rect 16028 20408 16080 20417
rect 16304 20408 16356 20460
rect 12440 20315 12492 20324
rect 12440 20281 12449 20315
rect 12449 20281 12483 20315
rect 12483 20281 12492 20315
rect 12440 20272 12492 20281
rect 5632 20204 5684 20256
rect 8300 20204 8352 20256
rect 8944 20204 8996 20256
rect 12532 20247 12584 20256
rect 12532 20213 12541 20247
rect 12541 20213 12575 20247
rect 12575 20213 12584 20247
rect 12532 20204 12584 20213
rect 15384 20340 15436 20392
rect 13452 20204 13504 20256
rect 14372 20204 14424 20256
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 6828 20043 6880 20052
rect 6828 20009 6837 20043
rect 6837 20009 6871 20043
rect 6871 20009 6880 20043
rect 6828 20000 6880 20009
rect 13176 20000 13228 20052
rect 13820 19975 13872 19984
rect 13820 19941 13829 19975
rect 13829 19941 13863 19975
rect 13863 19941 13872 19975
rect 13820 19932 13872 19941
rect 14464 20000 14516 20052
rect 16304 20000 16356 20052
rect 14832 19932 14884 19984
rect 5356 19864 5408 19916
rect 13452 19864 13504 19916
rect 6184 19796 6236 19848
rect 6736 19796 6788 19848
rect 8944 19796 8996 19848
rect 12532 19796 12584 19848
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 14740 19864 14792 19916
rect 15384 19796 15436 19848
rect 28540 19839 28592 19848
rect 28540 19805 28549 19839
rect 28549 19805 28583 19839
rect 28583 19805 28592 19839
rect 28540 19796 28592 19805
rect 6368 19728 6420 19780
rect 15660 19728 15712 19780
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 16764 19703 16816 19712
rect 16764 19669 16773 19703
rect 16773 19669 16807 19703
rect 16807 19669 16816 19703
rect 16764 19660 16816 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 6184 19499 6236 19508
rect 6184 19465 6193 19499
rect 6193 19465 6227 19499
rect 6227 19465 6236 19499
rect 6184 19456 6236 19465
rect 6368 19499 6420 19508
rect 6368 19465 6377 19499
rect 6377 19465 6411 19499
rect 6411 19465 6420 19499
rect 6368 19456 6420 19465
rect 7380 19499 7432 19508
rect 7380 19465 7389 19499
rect 7389 19465 7423 19499
rect 7423 19465 7432 19499
rect 7380 19456 7432 19465
rect 15660 19499 15712 19508
rect 15660 19465 15669 19499
rect 15669 19465 15703 19499
rect 15703 19465 15712 19499
rect 15660 19456 15712 19465
rect 5356 19388 5408 19440
rect 8852 19320 8904 19372
rect 15844 19363 15896 19372
rect 15844 19329 15853 19363
rect 15853 19329 15887 19363
rect 15887 19329 15896 19363
rect 15844 19320 15896 19329
rect 16764 19388 16816 19440
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 16672 19320 16724 19372
rect 17960 19320 18012 19372
rect 6920 19252 6972 19304
rect 7196 19295 7248 19304
rect 7196 19261 7205 19295
rect 7205 19261 7239 19295
rect 7239 19261 7248 19295
rect 7196 19252 7248 19261
rect 9772 19252 9824 19304
rect 8760 19116 8812 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 7012 18912 7064 18964
rect 22100 18844 22152 18896
rect 5356 18819 5408 18828
rect 5356 18785 5365 18819
rect 5365 18785 5399 18819
rect 5399 18785 5408 18819
rect 5356 18776 5408 18785
rect 8944 18819 8996 18828
rect 8944 18785 8953 18819
rect 8953 18785 8987 18819
rect 8987 18785 8996 18819
rect 8944 18776 8996 18785
rect 21088 18776 21140 18828
rect 5632 18751 5684 18760
rect 5632 18717 5666 18751
rect 5666 18717 5684 18751
rect 5632 18708 5684 18717
rect 19248 18708 19300 18760
rect 20904 18708 20956 18760
rect 21180 18751 21232 18760
rect 21180 18717 21189 18751
rect 21189 18717 21223 18751
rect 21223 18717 21232 18751
rect 21180 18708 21232 18717
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 22100 18708 22152 18760
rect 9036 18640 9088 18692
rect 19616 18640 19668 18692
rect 20720 18640 20772 18692
rect 23664 18640 23716 18692
rect 23940 18751 23992 18760
rect 23940 18717 23949 18751
rect 23949 18717 23983 18751
rect 23983 18717 23992 18751
rect 23940 18708 23992 18717
rect 25504 18640 25556 18692
rect 27528 18640 27580 18692
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 21088 18572 21140 18624
rect 23112 18572 23164 18624
rect 23480 18572 23532 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 23664 18368 23716 18420
rect 8760 18275 8812 18284
rect 8760 18241 8769 18275
rect 8769 18241 8803 18275
rect 8803 18241 8812 18275
rect 8760 18232 8812 18241
rect 8852 18275 8904 18284
rect 8852 18241 8881 18275
rect 8881 18241 8904 18275
rect 13176 18300 13228 18352
rect 8852 18232 8904 18241
rect 9864 18232 9916 18284
rect 11336 18164 11388 18216
rect 16120 18232 16172 18284
rect 17960 18275 18012 18284
rect 17960 18241 17969 18275
rect 17969 18241 18003 18275
rect 18003 18241 18012 18275
rect 17960 18232 18012 18241
rect 18696 18232 18748 18284
rect 19248 18232 19300 18284
rect 20444 18275 20496 18284
rect 20444 18241 20478 18275
rect 20478 18241 20496 18275
rect 20444 18232 20496 18241
rect 22284 18275 22336 18284
rect 22284 18241 22318 18275
rect 22318 18241 22336 18275
rect 22284 18232 22336 18241
rect 23756 18275 23808 18284
rect 23756 18241 23790 18275
rect 23790 18241 23808 18275
rect 23756 18232 23808 18241
rect 15936 18164 15988 18216
rect 18512 18164 18564 18216
rect 25228 18275 25280 18284
rect 25228 18241 25262 18275
rect 25262 18241 25280 18275
rect 25228 18232 25280 18241
rect 9772 18028 9824 18080
rect 10508 18028 10560 18080
rect 15200 18071 15252 18080
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 18328 18028 18380 18080
rect 19248 18071 19300 18080
rect 19248 18037 19257 18071
rect 19257 18037 19291 18071
rect 19291 18037 19300 18071
rect 19248 18028 19300 18037
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 24860 18071 24912 18080
rect 24860 18037 24869 18071
rect 24869 18037 24903 18071
rect 24903 18037 24912 18071
rect 24860 18028 24912 18037
rect 26240 18028 26292 18080
rect 26516 18028 26568 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 16120 17824 16172 17876
rect 19616 17867 19668 17876
rect 19616 17833 19625 17867
rect 19625 17833 19659 17867
rect 19659 17833 19668 17867
rect 19616 17824 19668 17833
rect 22284 17824 22336 17876
rect 23940 17824 23992 17876
rect 24032 17867 24084 17876
rect 24032 17833 24041 17867
rect 24041 17833 24075 17867
rect 24075 17833 24084 17867
rect 24032 17824 24084 17833
rect 25228 17824 25280 17876
rect 10232 17620 10284 17672
rect 10784 17620 10836 17672
rect 14740 17620 14792 17672
rect 18328 17620 18380 17672
rect 18420 17620 18472 17672
rect 21180 17756 21232 17808
rect 21456 17756 21508 17808
rect 18880 17620 18932 17672
rect 20812 17688 20864 17740
rect 21548 17688 21600 17740
rect 15200 17552 15252 17604
rect 18512 17595 18564 17604
rect 18512 17561 18521 17595
rect 18521 17561 18555 17595
rect 18555 17561 18564 17595
rect 20168 17663 20220 17672
rect 20168 17629 20177 17663
rect 20177 17629 20211 17663
rect 20211 17629 20220 17663
rect 20168 17620 20220 17629
rect 20904 17620 20956 17672
rect 21088 17663 21140 17672
rect 21088 17629 21097 17663
rect 21097 17629 21131 17663
rect 21131 17629 21140 17663
rect 21088 17620 21140 17629
rect 22560 17663 22612 17672
rect 22560 17629 22569 17663
rect 22569 17629 22603 17663
rect 22603 17629 22612 17663
rect 22560 17620 22612 17629
rect 18512 17552 18564 17561
rect 9864 17484 9916 17536
rect 18788 17527 18840 17536
rect 18788 17493 18797 17527
rect 18797 17493 18831 17527
rect 18831 17493 18840 17527
rect 18788 17484 18840 17493
rect 20168 17484 20220 17536
rect 22100 17552 22152 17604
rect 24768 17756 24820 17808
rect 23664 17731 23716 17740
rect 23664 17697 23673 17731
rect 23673 17697 23707 17731
rect 23707 17697 23716 17731
rect 23664 17688 23716 17697
rect 24032 17688 24084 17740
rect 25872 17688 25924 17740
rect 24308 17552 24360 17604
rect 24860 17552 24912 17604
rect 25412 17620 25464 17672
rect 26516 17663 26568 17672
rect 26516 17629 26525 17663
rect 26525 17629 26559 17663
rect 26559 17629 26568 17663
rect 26516 17620 26568 17629
rect 20996 17484 21048 17536
rect 24400 17527 24452 17536
rect 24400 17493 24409 17527
rect 24409 17493 24443 17527
rect 24443 17493 24452 17527
rect 24400 17484 24452 17493
rect 25596 17484 25648 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 20444 17280 20496 17332
rect 21180 17280 21232 17332
rect 21456 17323 21508 17332
rect 21456 17289 21465 17323
rect 21465 17289 21499 17323
rect 21499 17289 21508 17323
rect 21456 17280 21508 17289
rect 22560 17280 22612 17332
rect 23756 17280 23808 17332
rect 25596 17323 25648 17332
rect 25596 17289 25605 17323
rect 25605 17289 25639 17323
rect 25639 17289 25648 17323
rect 25596 17280 25648 17289
rect 10232 17212 10284 17264
rect 11520 17212 11572 17264
rect 18788 17212 18840 17264
rect 20812 17212 20864 17264
rect 11244 17144 11296 17196
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 20720 17187 20772 17196
rect 20720 17153 20729 17187
rect 20729 17153 20763 17187
rect 20763 17153 20772 17187
rect 20720 17144 20772 17153
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 20996 17187 21048 17196
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 20996 17144 21048 17153
rect 22100 17144 22152 17196
rect 23112 17187 23164 17196
rect 23112 17153 23121 17187
rect 23121 17153 23155 17187
rect 23155 17153 23164 17187
rect 23112 17144 23164 17153
rect 24400 17212 24452 17264
rect 24768 17212 24820 17264
rect 23480 17187 23532 17196
rect 23480 17153 23489 17187
rect 23489 17153 23523 17187
rect 23523 17153 23532 17187
rect 23480 17144 23532 17153
rect 25504 17144 25556 17196
rect 18144 17076 18196 17128
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 19708 17051 19760 17060
rect 19708 17017 19717 17051
rect 19717 17017 19751 17051
rect 19751 17017 19760 17051
rect 19708 17008 19760 17017
rect 25412 17051 25464 17060
rect 25412 17017 25421 17051
rect 25421 17017 25455 17051
rect 25455 17017 25464 17051
rect 25412 17008 25464 17017
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 11152 16940 11204 16992
rect 12164 16940 12216 16992
rect 16856 16940 16908 16992
rect 19800 16983 19852 16992
rect 19800 16949 19809 16983
rect 19809 16949 19843 16983
rect 19843 16949 19852 16983
rect 19800 16940 19852 16949
rect 20628 16940 20680 16992
rect 21088 16940 21140 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 9956 16668 10008 16720
rect 10784 16711 10836 16720
rect 10784 16677 10793 16711
rect 10793 16677 10827 16711
rect 10827 16677 10836 16711
rect 10784 16668 10836 16677
rect 11244 16736 11296 16788
rect 12164 16779 12216 16788
rect 12164 16745 12173 16779
rect 12173 16745 12207 16779
rect 12207 16745 12216 16779
rect 12164 16736 12216 16745
rect 5540 16532 5592 16584
rect 7656 16532 7708 16584
rect 8300 16532 8352 16584
rect 9864 16575 9916 16584
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 9956 16575 10008 16584
rect 9956 16541 9965 16575
rect 9965 16541 9999 16575
rect 9999 16541 10008 16575
rect 9956 16532 10008 16541
rect 11152 16600 11204 16652
rect 11612 16668 11664 16720
rect 11520 16600 11572 16652
rect 18328 16736 18380 16788
rect 18420 16779 18472 16788
rect 18420 16745 18429 16779
rect 18429 16745 18463 16779
rect 18463 16745 18472 16779
rect 18420 16736 18472 16745
rect 19708 16736 19760 16788
rect 25596 16779 25648 16788
rect 25596 16745 25605 16779
rect 25605 16745 25639 16779
rect 25639 16745 25648 16779
rect 25596 16736 25648 16745
rect 18880 16711 18932 16720
rect 18880 16677 18889 16711
rect 18889 16677 18923 16711
rect 18923 16677 18932 16711
rect 18880 16668 18932 16677
rect 26240 16600 26292 16652
rect 11060 16507 11112 16516
rect 11060 16473 11069 16507
rect 11069 16473 11103 16507
rect 11103 16473 11112 16507
rect 11060 16464 11112 16473
rect 11152 16507 11204 16516
rect 11152 16473 11161 16507
rect 11161 16473 11195 16507
rect 11195 16473 11204 16507
rect 12532 16575 12584 16584
rect 12532 16541 12541 16575
rect 12541 16541 12575 16575
rect 12575 16541 12584 16575
rect 12532 16532 12584 16541
rect 16856 16575 16908 16584
rect 16856 16541 16890 16575
rect 16890 16541 16908 16575
rect 16856 16532 16908 16541
rect 17316 16532 17368 16584
rect 19800 16532 19852 16584
rect 25504 16575 25556 16584
rect 25504 16541 25513 16575
rect 25513 16541 25547 16575
rect 25547 16541 25556 16575
rect 25504 16532 25556 16541
rect 25872 16575 25924 16584
rect 25872 16541 25881 16575
rect 25881 16541 25915 16575
rect 25915 16541 25924 16575
rect 25872 16532 25924 16541
rect 11152 16464 11204 16473
rect 5816 16396 5868 16448
rect 6276 16396 6328 16448
rect 7656 16396 7708 16448
rect 11520 16396 11572 16448
rect 18236 16439 18288 16448
rect 18236 16405 18245 16439
rect 18245 16405 18279 16439
rect 18279 16405 18288 16439
rect 18236 16396 18288 16405
rect 18512 16507 18564 16516
rect 18512 16473 18521 16507
rect 18521 16473 18555 16507
rect 18555 16473 18564 16507
rect 18512 16464 18564 16473
rect 24860 16396 24912 16448
rect 25596 16396 25648 16448
rect 28264 16439 28316 16448
rect 28264 16405 28273 16439
rect 28273 16405 28307 16439
rect 28307 16405 28316 16439
rect 28264 16396 28316 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 5540 16235 5592 16244
rect 5540 16201 5549 16235
rect 5549 16201 5583 16235
rect 5583 16201 5592 16235
rect 5540 16192 5592 16201
rect 8300 16192 8352 16244
rect 8576 16192 8628 16244
rect 9956 16192 10008 16244
rect 11152 16192 11204 16244
rect 18236 16192 18288 16244
rect 18512 16192 18564 16244
rect 25504 16192 25556 16244
rect 28448 16235 28500 16244
rect 28448 16201 28457 16235
rect 28457 16201 28491 16235
rect 28491 16201 28500 16235
rect 28448 16192 28500 16201
rect 848 16056 900 16108
rect 3424 15988 3476 16040
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 6000 16099 6052 16108
rect 6000 16065 6009 16099
rect 6009 16065 6043 16099
rect 6043 16065 6052 16099
rect 6000 16056 6052 16065
rect 9496 16124 9548 16176
rect 12164 16124 12216 16176
rect 18144 16124 18196 16176
rect 21456 16124 21508 16176
rect 3240 15852 3292 15904
rect 8300 16056 8352 16108
rect 10324 16099 10376 16108
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 10600 16056 10652 16108
rect 17776 16099 17828 16108
rect 17776 16065 17794 16099
rect 17794 16065 17828 16099
rect 17776 16056 17828 16065
rect 18328 16056 18380 16108
rect 10692 16031 10744 16040
rect 10692 15997 10701 16031
rect 10701 15997 10735 16031
rect 10735 15997 10744 16031
rect 10692 15988 10744 15997
rect 12072 16031 12124 16040
rect 12072 15997 12081 16031
rect 12081 15997 12115 16031
rect 12115 15997 12124 16031
rect 12072 15988 12124 15997
rect 8484 15920 8536 15972
rect 7288 15852 7340 15904
rect 9036 15852 9088 15904
rect 13728 15852 13780 15904
rect 17316 15852 17368 15904
rect 23296 16099 23348 16108
rect 23296 16065 23305 16099
rect 23305 16065 23339 16099
rect 23339 16065 23348 16099
rect 23296 16056 23348 16065
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 22192 15988 22244 16040
rect 23388 15988 23440 16040
rect 24308 16056 24360 16108
rect 24860 16056 24912 16108
rect 28264 16099 28316 16108
rect 28264 16065 28273 16099
rect 28273 16065 28307 16099
rect 28307 16065 28316 16099
rect 28264 16056 28316 16065
rect 18144 15895 18196 15904
rect 18144 15861 18153 15895
rect 18153 15861 18187 15895
rect 18187 15861 18196 15895
rect 18144 15852 18196 15861
rect 19156 15895 19208 15904
rect 19156 15861 19165 15895
rect 19165 15861 19199 15895
rect 19199 15861 19208 15895
rect 19156 15852 19208 15861
rect 26516 15920 26568 15972
rect 25228 15852 25280 15904
rect 28172 15895 28224 15904
rect 28172 15861 28181 15895
rect 28181 15861 28215 15895
rect 28215 15861 28224 15895
rect 28172 15852 28224 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 3424 15691 3476 15700
rect 3424 15657 3433 15691
rect 3433 15657 3467 15691
rect 3467 15657 3476 15691
rect 3424 15648 3476 15657
rect 7656 15648 7708 15700
rect 11060 15691 11112 15700
rect 11060 15657 11069 15691
rect 11069 15657 11103 15691
rect 11103 15657 11112 15691
rect 11060 15648 11112 15657
rect 8024 15580 8076 15632
rect 11612 15648 11664 15700
rect 12532 15648 12584 15700
rect 17776 15648 17828 15700
rect 18144 15691 18196 15700
rect 18144 15657 18153 15691
rect 18153 15657 18187 15691
rect 18187 15657 18196 15691
rect 18144 15648 18196 15657
rect 3240 15487 3292 15496
rect 3240 15453 3249 15487
rect 3249 15453 3283 15487
rect 3283 15453 3292 15487
rect 3240 15444 3292 15453
rect 6276 15555 6328 15564
rect 6276 15521 6285 15555
rect 6285 15521 6319 15555
rect 6319 15521 6328 15555
rect 6276 15512 6328 15521
rect 8484 15555 8536 15564
rect 8484 15521 8493 15555
rect 8493 15521 8527 15555
rect 8527 15521 8536 15555
rect 8484 15512 8536 15521
rect 6000 15444 6052 15496
rect 7288 15444 7340 15496
rect 8300 15419 8352 15428
rect 7840 15308 7892 15360
rect 8024 15308 8076 15360
rect 8300 15385 8309 15419
rect 8309 15385 8343 15419
rect 8343 15385 8352 15419
rect 8300 15376 8352 15385
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 10968 15444 11020 15496
rect 9036 15376 9088 15428
rect 11336 15444 11388 15496
rect 11520 15487 11572 15496
rect 11520 15453 11554 15487
rect 11554 15453 11572 15487
rect 11520 15444 11572 15453
rect 19156 15512 19208 15564
rect 18236 15487 18288 15496
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 19892 15487 19944 15496
rect 19892 15453 19901 15487
rect 19901 15453 19935 15487
rect 19935 15453 19944 15487
rect 19892 15444 19944 15453
rect 19984 15487 20036 15496
rect 19984 15453 19994 15487
rect 19994 15453 20028 15487
rect 20028 15453 20036 15487
rect 19984 15444 20036 15453
rect 19340 15376 19392 15428
rect 20260 15419 20312 15428
rect 20260 15385 20269 15419
rect 20269 15385 20303 15419
rect 20303 15385 20312 15419
rect 20260 15376 20312 15385
rect 10508 15308 10560 15360
rect 19432 15308 19484 15360
rect 20628 15444 20680 15496
rect 20812 15444 20864 15496
rect 21548 15487 21600 15496
rect 21548 15453 21558 15487
rect 21558 15453 21592 15487
rect 21592 15453 21600 15487
rect 21548 15444 21600 15453
rect 21732 15308 21784 15360
rect 22100 15308 22152 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 8484 15104 8536 15156
rect 10692 15104 10744 15156
rect 10968 15147 11020 15156
rect 10968 15113 10977 15147
rect 10977 15113 11011 15147
rect 11011 15113 11020 15147
rect 10968 15104 11020 15113
rect 7564 15011 7616 15020
rect 7564 14977 7598 15011
rect 7598 14977 7616 15011
rect 7564 14968 7616 14977
rect 10508 15079 10560 15088
rect 10508 15045 10517 15079
rect 10517 15045 10551 15079
rect 10551 15045 10560 15079
rect 10508 15036 10560 15045
rect 13728 15036 13780 15088
rect 9680 14968 9732 15020
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 12532 14968 12584 15020
rect 13452 15011 13504 15020
rect 13452 14977 13461 15011
rect 13461 14977 13495 15011
rect 13495 14977 13504 15011
rect 13452 14968 13504 14977
rect 13636 14968 13688 15020
rect 23296 15104 23348 15156
rect 17224 15036 17276 15088
rect 22100 15079 22152 15088
rect 22100 15045 22109 15079
rect 22109 15045 22143 15079
rect 22143 15045 22152 15079
rect 22100 15036 22152 15045
rect 22192 15079 22244 15088
rect 22192 15045 22201 15079
rect 22201 15045 22235 15079
rect 22235 15045 22244 15079
rect 22192 15036 22244 15045
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 10600 14943 10652 14952
rect 10600 14909 10609 14943
rect 10609 14909 10643 14943
rect 10643 14909 10652 14943
rect 10600 14900 10652 14909
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 14924 15011 14976 15020
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 17316 14968 17368 15020
rect 21732 14968 21784 15020
rect 23480 14968 23532 15020
rect 10324 14764 10376 14816
rect 16212 14764 16264 14816
rect 18328 14764 18380 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 7564 14560 7616 14612
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 13728 14560 13780 14612
rect 19340 14560 19392 14612
rect 19984 14560 20036 14612
rect 13360 14492 13412 14544
rect 13636 14492 13688 14544
rect 8484 14424 8536 14476
rect 7840 14399 7892 14408
rect 7840 14365 7849 14399
rect 7849 14365 7883 14399
rect 7883 14365 7892 14399
rect 7840 14356 7892 14365
rect 8300 14356 8352 14408
rect 9772 14356 9824 14408
rect 10232 14356 10284 14408
rect 13452 14399 13504 14408
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 14924 14492 14976 14544
rect 13360 14288 13412 14340
rect 13636 14331 13688 14340
rect 13636 14297 13645 14331
rect 13645 14297 13679 14331
rect 13679 14297 13688 14331
rect 13636 14288 13688 14297
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 18236 14424 18288 14476
rect 17224 14399 17276 14408
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 18328 14399 18380 14408
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 18420 14356 18472 14408
rect 19708 14492 19760 14544
rect 19892 14492 19944 14544
rect 20812 14535 20864 14544
rect 20812 14501 20821 14535
rect 20821 14501 20855 14535
rect 20855 14501 20864 14535
rect 20812 14492 20864 14501
rect 19340 14467 19392 14476
rect 19340 14433 19349 14467
rect 19349 14433 19383 14467
rect 19383 14433 19392 14467
rect 19340 14424 19392 14433
rect 13452 14220 13504 14272
rect 15476 14288 15528 14340
rect 18880 14356 18932 14408
rect 20260 14424 20312 14476
rect 19708 14356 19760 14408
rect 21548 14288 21600 14340
rect 15292 14220 15344 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 25596 14059 25648 14068
rect 25596 14025 25605 14059
rect 25605 14025 25639 14059
rect 25639 14025 25648 14059
rect 25596 14016 25648 14025
rect 18696 13991 18748 14000
rect 18696 13957 18705 13991
rect 18705 13957 18739 13991
rect 18739 13957 18748 13991
rect 18696 13948 18748 13957
rect 16212 13880 16264 13932
rect 25320 13923 25372 13932
rect 25320 13889 25329 13923
rect 25329 13889 25363 13923
rect 25363 13889 25372 13923
rect 25320 13880 25372 13889
rect 25688 13923 25740 13932
rect 25688 13889 25697 13923
rect 25697 13889 25731 13923
rect 25731 13889 25740 13923
rect 25688 13880 25740 13889
rect 25412 13812 25464 13864
rect 17224 13719 17276 13728
rect 17224 13685 17233 13719
rect 17233 13685 17267 13719
rect 17267 13685 17276 13719
rect 17224 13676 17276 13685
rect 24860 13719 24912 13728
rect 24860 13685 24869 13719
rect 24869 13685 24903 13719
rect 24903 13685 24912 13719
rect 24860 13676 24912 13685
rect 25044 13719 25096 13728
rect 25044 13685 25053 13719
rect 25053 13685 25087 13719
rect 25087 13685 25096 13719
rect 25044 13676 25096 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 13360 13472 13412 13524
rect 15476 13472 15528 13524
rect 25044 13472 25096 13524
rect 25688 13472 25740 13524
rect 12072 13336 12124 13388
rect 16764 13336 16816 13388
rect 21824 13336 21876 13388
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 12624 13243 12676 13252
rect 12624 13209 12658 13243
rect 12658 13209 12676 13243
rect 12624 13200 12676 13209
rect 17224 13268 17276 13320
rect 20720 13268 20772 13320
rect 21456 13268 21508 13320
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 24492 13311 24544 13320
rect 24492 13277 24501 13311
rect 24501 13277 24535 13311
rect 24535 13277 24544 13311
rect 24492 13268 24544 13277
rect 16580 13200 16632 13252
rect 17040 13200 17092 13252
rect 24860 13268 24912 13320
rect 15476 13132 15528 13184
rect 16028 13175 16080 13184
rect 16028 13141 16037 13175
rect 16037 13141 16071 13175
rect 16071 13141 16080 13175
rect 16028 13132 16080 13141
rect 16120 13175 16172 13184
rect 16120 13141 16129 13175
rect 16129 13141 16163 13175
rect 16163 13141 16172 13175
rect 16120 13132 16172 13141
rect 22008 13132 22060 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 16028 12860 16080 12912
rect 16120 12792 16172 12844
rect 21824 12835 21876 12844
rect 21824 12801 21833 12835
rect 21833 12801 21867 12835
rect 21867 12801 21876 12835
rect 21824 12792 21876 12801
rect 22008 12860 22060 12912
rect 22376 12792 22428 12844
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 25320 12928 25372 12980
rect 25596 12928 25648 12980
rect 23296 12835 23348 12844
rect 23296 12801 23305 12835
rect 23305 12801 23339 12835
rect 23339 12801 23348 12835
rect 23296 12792 23348 12801
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 16948 12767 17000 12776
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 21364 12767 21416 12776
rect 21364 12733 21373 12767
rect 21373 12733 21407 12767
rect 21407 12733 21416 12767
rect 21364 12724 21416 12733
rect 24860 12724 24912 12776
rect 17960 12656 18012 12708
rect 21640 12699 21692 12708
rect 21640 12665 21649 12699
rect 21649 12665 21683 12699
rect 21683 12665 21692 12699
rect 21640 12656 21692 12665
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 11520 12384 11572 12436
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 16948 12384 17000 12436
rect 21732 12384 21784 12436
rect 22376 12384 22428 12436
rect 23388 12384 23440 12436
rect 21548 12316 21600 12368
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 11704 12180 11756 12232
rect 21456 12291 21508 12300
rect 21456 12257 21465 12291
rect 21465 12257 21499 12291
rect 21499 12257 21508 12291
rect 21456 12248 21508 12257
rect 13452 12180 13504 12232
rect 15200 12180 15252 12232
rect 21640 12180 21692 12232
rect 22284 12180 22336 12232
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 23296 12291 23348 12300
rect 23296 12257 23305 12291
rect 23305 12257 23339 12291
rect 23339 12257 23348 12291
rect 23296 12248 23348 12257
rect 24492 12180 24544 12232
rect 9588 12087 9640 12096
rect 9588 12053 9597 12087
rect 9597 12053 9631 12087
rect 9631 12053 9640 12087
rect 9588 12044 9640 12053
rect 22376 12087 22428 12096
rect 22376 12053 22385 12087
rect 22385 12053 22419 12087
rect 22419 12053 22428 12087
rect 22376 12044 22428 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 16580 11840 16632 11892
rect 9588 11772 9640 11824
rect 16120 11772 16172 11824
rect 16212 11815 16264 11824
rect 16212 11781 16221 11815
rect 16221 11781 16255 11815
rect 16255 11781 16264 11815
rect 16212 11772 16264 11781
rect 16764 11815 16816 11824
rect 16764 11781 16773 11815
rect 16773 11781 16807 11815
rect 16807 11781 16816 11815
rect 16764 11772 16816 11781
rect 21180 11772 21232 11824
rect 23020 11772 23072 11824
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 9036 11636 9088 11688
rect 16488 11636 16540 11688
rect 18788 11636 18840 11688
rect 16028 11611 16080 11620
rect 16028 11577 16037 11611
rect 16037 11577 16071 11611
rect 16071 11577 16080 11611
rect 16028 11568 16080 11577
rect 18052 11611 18104 11620
rect 18052 11577 18061 11611
rect 18061 11577 18095 11611
rect 18095 11577 18104 11611
rect 18052 11568 18104 11577
rect 10508 11543 10560 11552
rect 10508 11509 10517 11543
rect 10517 11509 10551 11543
rect 10551 11509 10560 11543
rect 10508 11500 10560 11509
rect 11336 11500 11388 11552
rect 15108 11500 15160 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 11704 11339 11756 11348
rect 11704 11305 11713 11339
rect 11713 11305 11747 11339
rect 11747 11305 11756 11339
rect 11704 11296 11756 11305
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 15476 11296 15528 11348
rect 21456 11296 21508 11348
rect 12072 11203 12124 11212
rect 12072 11169 12081 11203
rect 12081 11169 12115 11203
rect 12115 11169 12124 11203
rect 12072 11160 12124 11169
rect 15108 11203 15160 11212
rect 15108 11169 15117 11203
rect 15117 11169 15151 11203
rect 15151 11169 15160 11203
rect 15108 11160 15160 11169
rect 16028 11203 16080 11212
rect 16028 11169 16037 11203
rect 16037 11169 16071 11203
rect 16071 11169 16080 11203
rect 16028 11160 16080 11169
rect 9036 11092 9088 11144
rect 15200 11092 15252 11144
rect 16580 11228 16632 11280
rect 21640 11228 21692 11280
rect 21272 11160 21324 11212
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 9220 11067 9272 11076
rect 9220 11033 9254 11067
rect 9254 11033 9272 11067
rect 9220 11024 9272 11033
rect 9312 11024 9364 11076
rect 12900 11024 12952 11076
rect 15752 11024 15804 11076
rect 21364 11092 21416 11144
rect 21916 11160 21968 11212
rect 24492 11160 24544 11212
rect 22284 11135 22336 11144
rect 22284 11101 22293 11135
rect 22293 11101 22327 11135
rect 22327 11101 22336 11135
rect 22284 11092 22336 11101
rect 21548 11024 21600 11076
rect 22008 11024 22060 11076
rect 15476 10999 15528 11008
rect 15476 10965 15485 10999
rect 15485 10965 15519 10999
rect 15519 10965 15528 10999
rect 15476 10956 15528 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 9220 10752 9272 10804
rect 11704 10752 11756 10804
rect 9772 10684 9824 10736
rect 10140 10684 10192 10736
rect 12900 10795 12952 10804
rect 12900 10761 12909 10795
rect 12909 10761 12943 10795
rect 12943 10761 12952 10795
rect 12900 10752 12952 10761
rect 13176 10795 13228 10804
rect 13176 10761 13185 10795
rect 13185 10761 13219 10795
rect 13219 10761 13228 10795
rect 13176 10752 13228 10761
rect 15752 10752 15804 10804
rect 11336 10659 11388 10668
rect 11336 10625 11345 10659
rect 11345 10625 11379 10659
rect 11379 10625 11388 10659
rect 11336 10616 11388 10625
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 12716 10684 12768 10736
rect 14556 10684 14608 10736
rect 19524 10752 19576 10804
rect 21272 10752 21324 10804
rect 25596 10752 25648 10804
rect 19616 10684 19668 10736
rect 25136 10684 25188 10736
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 15200 10616 15252 10668
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 17960 10616 18012 10625
rect 18236 10616 18288 10668
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 8760 10591 8812 10600
rect 8760 10557 8769 10591
rect 8769 10557 8803 10591
rect 8803 10557 8812 10591
rect 8760 10548 8812 10557
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 18144 10548 18196 10600
rect 18788 10591 18840 10600
rect 18788 10557 18797 10591
rect 18797 10557 18831 10591
rect 18831 10557 18840 10591
rect 18788 10548 18840 10557
rect 19432 10591 19484 10600
rect 19432 10557 19441 10591
rect 19441 10557 19475 10591
rect 19475 10557 19484 10591
rect 19432 10548 19484 10557
rect 19524 10591 19576 10600
rect 19524 10557 19533 10591
rect 19533 10557 19567 10591
rect 19567 10557 19576 10591
rect 19524 10548 19576 10557
rect 24492 10659 24544 10668
rect 24492 10625 24501 10659
rect 24501 10625 24535 10659
rect 24535 10625 24544 10659
rect 24492 10616 24544 10625
rect 24768 10659 24820 10668
rect 24768 10625 24777 10659
rect 24777 10625 24811 10659
rect 24811 10625 24820 10659
rect 24768 10616 24820 10625
rect 24860 10616 24912 10668
rect 25964 10616 26016 10668
rect 19340 10480 19392 10532
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 18420 10412 18472 10464
rect 18788 10412 18840 10464
rect 19156 10412 19208 10464
rect 21364 10412 21416 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 10140 10251 10192 10260
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 11060 10208 11112 10260
rect 11888 10208 11940 10260
rect 15200 10251 15252 10260
rect 15200 10217 15209 10251
rect 15209 10217 15243 10251
rect 15243 10217 15252 10251
rect 15200 10208 15252 10217
rect 24768 10208 24820 10260
rect 940 10004 992 10056
rect 10784 10072 10836 10124
rect 11520 10072 11572 10124
rect 18420 10115 18472 10124
rect 18420 10081 18429 10115
rect 18429 10081 18463 10115
rect 18463 10081 18472 10115
rect 18420 10072 18472 10081
rect 18512 10115 18564 10124
rect 18512 10081 18521 10115
rect 18521 10081 18555 10115
rect 18555 10081 18564 10115
rect 18512 10072 18564 10081
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 12072 10004 12124 10056
rect 14464 10004 14516 10056
rect 15016 10047 15068 10056
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 15476 10004 15528 10056
rect 18144 10004 18196 10056
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 21364 10140 21416 10192
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 19064 10004 19116 10056
rect 24860 10140 24912 10192
rect 25136 10183 25188 10192
rect 25136 10149 25145 10183
rect 25145 10149 25179 10183
rect 25179 10149 25188 10183
rect 25136 10140 25188 10149
rect 24492 10115 24544 10124
rect 24492 10081 24501 10115
rect 24501 10081 24535 10115
rect 24535 10081 24544 10115
rect 24492 10072 24544 10081
rect 25596 10208 25648 10260
rect 26792 10208 26844 10260
rect 10600 9979 10652 9988
rect 10600 9945 10609 9979
rect 10609 9945 10643 9979
rect 10643 9945 10652 9979
rect 10600 9936 10652 9945
rect 10968 9936 11020 9988
rect 18604 9936 18656 9988
rect 19340 9936 19392 9988
rect 25964 10047 26016 10056
rect 25964 10013 25973 10047
rect 25973 10013 26007 10047
rect 26007 10013 26016 10047
rect 25964 10004 26016 10013
rect 28356 9936 28408 9988
rect 11060 9868 11112 9920
rect 11520 9868 11572 9920
rect 17960 9911 18012 9920
rect 17960 9877 17969 9911
rect 17969 9877 18003 9911
rect 18003 9877 18012 9911
rect 17960 9868 18012 9877
rect 18144 9868 18196 9920
rect 18512 9868 18564 9920
rect 19524 9868 19576 9920
rect 19708 9868 19760 9920
rect 24952 9911 25004 9920
rect 24952 9877 24961 9911
rect 24961 9877 24995 9911
rect 24995 9877 25004 9911
rect 24952 9868 25004 9877
rect 25228 9868 25280 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 10416 9664 10468 9716
rect 10692 9664 10744 9716
rect 11520 9707 11572 9716
rect 11520 9673 11529 9707
rect 11529 9673 11563 9707
rect 11563 9673 11572 9707
rect 11520 9664 11572 9673
rect 5816 9528 5868 9580
rect 9312 9596 9364 9648
rect 9956 9596 10008 9648
rect 14556 9639 14608 9648
rect 14556 9605 14565 9639
rect 14565 9605 14599 9639
rect 14599 9605 14608 9639
rect 14556 9596 14608 9605
rect 15016 9639 15068 9648
rect 15016 9605 15025 9639
rect 15025 9605 15059 9639
rect 15059 9605 15068 9639
rect 15016 9596 15068 9605
rect 15200 9639 15252 9648
rect 15200 9605 15209 9639
rect 15209 9605 15243 9639
rect 15243 9605 15252 9639
rect 15200 9596 15252 9605
rect 7288 9528 7340 9580
rect 9772 9528 9824 9580
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 12164 9528 12216 9580
rect 16028 9664 16080 9716
rect 18144 9664 18196 9716
rect 18236 9664 18288 9716
rect 19432 9707 19484 9716
rect 19432 9673 19441 9707
rect 19441 9673 19475 9707
rect 19475 9673 19484 9707
rect 19432 9664 19484 9673
rect 24952 9664 25004 9716
rect 19340 9596 19392 9648
rect 15384 9528 15436 9580
rect 18052 9528 18104 9580
rect 18604 9571 18656 9580
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 19064 9571 19116 9580
rect 19064 9537 19073 9571
rect 19073 9537 19107 9571
rect 19107 9537 19116 9571
rect 19064 9528 19116 9537
rect 19156 9528 19208 9580
rect 21548 9528 21600 9580
rect 22008 9571 22060 9580
rect 9404 9460 9456 9512
rect 14464 9460 14516 9512
rect 20076 9460 20128 9512
rect 21180 9503 21232 9512
rect 21180 9469 21189 9503
rect 21189 9469 21223 9503
rect 21223 9469 21232 9503
rect 21180 9460 21232 9469
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 25412 9639 25464 9648
rect 25412 9605 25421 9639
rect 25421 9605 25455 9639
rect 25455 9605 25464 9639
rect 25412 9596 25464 9605
rect 25596 9639 25648 9648
rect 25596 9605 25605 9639
rect 25605 9605 25639 9639
rect 25639 9605 25648 9639
rect 25596 9596 25648 9605
rect 21916 9503 21968 9512
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 24584 9528 24636 9580
rect 25228 9528 25280 9580
rect 8760 9392 8812 9444
rect 10784 9392 10836 9444
rect 20720 9392 20772 9444
rect 22008 9392 22060 9444
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 11152 9324 11204 9376
rect 14924 9324 14976 9376
rect 22468 9324 22520 9376
rect 23940 9367 23992 9376
rect 23940 9333 23949 9367
rect 23949 9333 23983 9367
rect 23983 9333 23992 9367
rect 23940 9324 23992 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 5816 9027 5868 9036
rect 5816 8993 5825 9027
rect 5825 8993 5859 9027
rect 5859 8993 5868 9027
rect 5816 8984 5868 8993
rect 10140 9052 10192 9104
rect 10600 9120 10652 9172
rect 12164 9163 12216 9172
rect 12164 9129 12173 9163
rect 12173 9129 12207 9163
rect 12207 9129 12216 9163
rect 12164 9120 12216 9129
rect 15292 9120 15344 9172
rect 19524 9052 19576 9104
rect 22376 9120 22428 9172
rect 25964 9120 26016 9172
rect 10600 9027 10652 9036
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 10968 8984 11020 9036
rect 9956 8959 10008 8968
rect 9956 8925 9965 8959
rect 9965 8925 9999 8959
rect 9999 8925 10008 8959
rect 9956 8916 10008 8925
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 19708 9027 19760 9036
rect 19708 8993 19717 9027
rect 19717 8993 19751 9027
rect 19751 8993 19760 9027
rect 19708 8984 19760 8993
rect 21916 9052 21968 9104
rect 21548 8984 21600 9036
rect 21824 8984 21876 9036
rect 5632 8848 5684 8900
rect 10416 8848 10468 8900
rect 14280 8916 14332 8968
rect 15016 8916 15068 8968
rect 12348 8891 12400 8900
rect 12348 8857 12357 8891
rect 12357 8857 12391 8891
rect 12391 8857 12400 8891
rect 12348 8848 12400 8857
rect 14740 8848 14792 8900
rect 17960 8916 18012 8968
rect 19616 8959 19668 8968
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 20076 8959 20128 8968
rect 20076 8925 20085 8959
rect 20085 8925 20119 8959
rect 20119 8925 20128 8959
rect 20076 8916 20128 8925
rect 21916 8959 21968 8968
rect 21916 8925 21925 8959
rect 21925 8925 21959 8959
rect 21959 8925 21968 8959
rect 21916 8916 21968 8925
rect 22468 8959 22520 8968
rect 22468 8925 22477 8959
rect 22477 8925 22511 8959
rect 22511 8925 22520 8959
rect 22468 8916 22520 8925
rect 23940 8916 23992 8968
rect 18696 8848 18748 8900
rect 22008 8848 22060 8900
rect 7564 8780 7616 8832
rect 17224 8780 17276 8832
rect 18880 8780 18932 8832
rect 22100 8823 22152 8832
rect 22100 8789 22109 8823
rect 22109 8789 22143 8823
rect 22143 8789 22152 8823
rect 22100 8780 22152 8789
rect 22376 8823 22428 8832
rect 22376 8789 22385 8823
rect 22385 8789 22419 8823
rect 22419 8789 22428 8823
rect 22376 8780 22428 8789
rect 24584 8780 24636 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 7288 8619 7340 8628
rect 7288 8585 7297 8619
rect 7297 8585 7331 8619
rect 7331 8585 7340 8619
rect 7288 8576 7340 8585
rect 9772 8576 9824 8628
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 7840 8508 7892 8560
rect 9864 8508 9916 8560
rect 10416 8576 10468 8628
rect 14740 8619 14792 8628
rect 14740 8585 14749 8619
rect 14749 8585 14783 8619
rect 14783 8585 14792 8619
rect 14740 8576 14792 8585
rect 19064 8576 19116 8628
rect 21548 8576 21600 8628
rect 28356 8619 28408 8628
rect 28356 8585 28365 8619
rect 28365 8585 28399 8619
rect 28399 8585 28408 8619
rect 28356 8576 28408 8585
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 13176 8508 13228 8560
rect 14464 8508 14516 8560
rect 10968 8483 11020 8492
rect 9312 8415 9364 8424
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 15292 8440 15344 8492
rect 22100 8551 22152 8560
rect 22100 8517 22134 8551
rect 22134 8517 22152 8551
rect 22100 8508 22152 8517
rect 17224 8483 17276 8492
rect 17224 8449 17258 8483
rect 17258 8449 17276 8483
rect 17224 8440 17276 8449
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 19248 8440 19300 8492
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 28540 8483 28592 8492
rect 28540 8449 28549 8483
rect 28549 8449 28583 8483
rect 28583 8449 28592 8483
rect 28540 8440 28592 8449
rect 12348 8372 12400 8424
rect 15384 8372 15436 8424
rect 20720 8372 20772 8424
rect 19340 8304 19392 8356
rect 10784 8279 10836 8288
rect 10784 8245 10793 8279
rect 10793 8245 10827 8279
rect 10827 8245 10836 8279
rect 10784 8236 10836 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 9956 8032 10008 8084
rect 20168 8032 20220 8084
rect 19248 7939 19300 7948
rect 19248 7905 19257 7939
rect 19257 7905 19291 7939
rect 19291 7905 19300 7939
rect 19248 7896 19300 7905
rect 9312 7828 9364 7880
rect 19340 7828 19392 7880
rect 10784 7760 10836 7812
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 5448 2635 5500 2644
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 27068 2388 27120 2440
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 6458 49314 6514 50000
rect 24490 49314 24546 50000
rect 6458 49286 6592 49314
rect 6458 49200 6514 49286
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 6564 47054 6592 49286
rect 24490 49286 24624 49314
rect 24490 49200 24546 49286
rect 7104 47184 7156 47190
rect 7104 47126 7156 47132
rect 6552 47048 6604 47054
rect 6552 46990 6604 46996
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 7116 45490 7144 47126
rect 24596 45554 24624 49286
rect 24504 45526 24624 45554
rect 7104 45484 7156 45490
rect 7104 45426 7156 45432
rect 12348 45484 12400 45490
rect 12348 45426 12400 45432
rect 8208 45416 8260 45422
rect 8208 45358 8260 45364
rect 12072 45416 12124 45422
rect 12072 45358 12124 45364
rect 7288 45280 7340 45286
rect 7288 45222 7340 45228
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 7300 44810 7328 45222
rect 7288 44804 7340 44810
rect 7288 44746 7340 44752
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 8220 41426 8248 45358
rect 12084 45082 12112 45358
rect 12256 45348 12308 45354
rect 12256 45290 12308 45296
rect 12164 45280 12216 45286
rect 12164 45222 12216 45228
rect 12072 45076 12124 45082
rect 12072 45018 12124 45024
rect 9588 44940 9640 44946
rect 9588 44882 9640 44888
rect 8944 44736 8996 44742
rect 8944 44678 8996 44684
rect 8956 44470 8984 44678
rect 8944 44464 8996 44470
rect 8944 44406 8996 44412
rect 9600 44402 9628 44882
rect 11520 44804 11572 44810
rect 11520 44746 11572 44752
rect 9588 44396 9640 44402
rect 9588 44338 9640 44344
rect 8576 44192 8628 44198
rect 8576 44134 8628 44140
rect 8588 43790 8616 44134
rect 9600 43994 9628 44338
rect 9772 44328 9824 44334
rect 9772 44270 9824 44276
rect 9784 44146 9812 44270
rect 9784 44118 9904 44146
rect 9876 43994 9904 44118
rect 11532 43994 11560 44746
rect 11888 44736 11940 44742
rect 11888 44678 11940 44684
rect 11704 44396 11756 44402
rect 11704 44338 11756 44344
rect 9588 43988 9640 43994
rect 9588 43930 9640 43936
rect 9864 43988 9916 43994
rect 9864 43930 9916 43936
rect 11520 43988 11572 43994
rect 11520 43930 11572 43936
rect 8576 43784 8628 43790
rect 8576 43726 8628 43732
rect 9600 42770 9628 43930
rect 11716 43790 11744 44338
rect 11796 44192 11848 44198
rect 11796 44134 11848 44140
rect 11704 43784 11756 43790
rect 11704 43726 11756 43732
rect 11716 43450 11744 43726
rect 11704 43444 11756 43450
rect 11704 43386 11756 43392
rect 11716 43314 11744 43386
rect 11808 43314 11836 44134
rect 11900 43858 11928 44678
rect 12084 44402 12112 45018
rect 12176 44810 12204 45222
rect 12268 44878 12296 45290
rect 12256 44872 12308 44878
rect 12256 44814 12308 44820
rect 12164 44804 12216 44810
rect 12164 44746 12216 44752
rect 12072 44396 12124 44402
rect 12072 44338 12124 44344
rect 11888 43852 11940 43858
rect 11888 43794 11940 43800
rect 12176 43654 12204 44746
rect 12268 44538 12296 44814
rect 12256 44532 12308 44538
rect 12256 44474 12308 44480
rect 12360 43858 12388 45426
rect 12440 45280 12492 45286
rect 12440 45222 12492 45228
rect 12452 43994 12480 45222
rect 12532 44940 12584 44946
rect 12532 44882 12584 44888
rect 13544 44940 13596 44946
rect 13544 44882 13596 44888
rect 12544 44470 12572 44882
rect 12624 44804 12676 44810
rect 12624 44746 12676 44752
rect 12532 44464 12584 44470
rect 12532 44406 12584 44412
rect 12440 43988 12492 43994
rect 12440 43930 12492 43936
rect 12348 43852 12400 43858
rect 12348 43794 12400 43800
rect 12164 43648 12216 43654
rect 12164 43590 12216 43596
rect 12544 43314 12572 44406
rect 12636 43790 12664 44746
rect 13268 44532 13320 44538
rect 13268 44474 13320 44480
rect 13176 44396 13228 44402
rect 13176 44338 13228 44344
rect 12716 44192 12768 44198
rect 12716 44134 12768 44140
rect 12728 43858 12756 44134
rect 13188 43994 13216 44338
rect 13280 43994 13308 44474
rect 13556 44402 13584 44882
rect 13820 44872 13872 44878
rect 13820 44814 13872 44820
rect 13544 44396 13596 44402
rect 13544 44338 13596 44344
rect 13176 43988 13228 43994
rect 13176 43930 13228 43936
rect 13268 43988 13320 43994
rect 13268 43930 13320 43936
rect 12992 43920 13044 43926
rect 12992 43862 13044 43868
rect 12716 43852 12768 43858
rect 12716 43794 12768 43800
rect 13004 43790 13032 43862
rect 13832 43790 13860 44814
rect 14464 44804 14516 44810
rect 14464 44746 14516 44752
rect 14476 44402 14504 44746
rect 14464 44396 14516 44402
rect 14464 44338 14516 44344
rect 12624 43784 12676 43790
rect 12624 43726 12676 43732
rect 12992 43784 13044 43790
rect 12992 43726 13044 43732
rect 13176 43784 13228 43790
rect 13176 43726 13228 43732
rect 13820 43784 13872 43790
rect 13820 43726 13872 43732
rect 14648 43784 14700 43790
rect 14648 43726 14700 43732
rect 12624 43648 12676 43654
rect 12624 43590 12676 43596
rect 12808 43648 12860 43654
rect 12808 43590 12860 43596
rect 11704 43308 11756 43314
rect 11704 43250 11756 43256
rect 11796 43308 11848 43314
rect 11796 43250 11848 43256
rect 12532 43308 12584 43314
rect 12532 43250 12584 43256
rect 12440 43240 12492 43246
rect 12440 43182 12492 43188
rect 11336 43104 11388 43110
rect 11336 43046 11388 43052
rect 9588 42764 9640 42770
rect 9588 42706 9640 42712
rect 8220 41398 8340 41426
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 7932 38956 7984 38962
rect 7932 38898 7984 38904
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 7944 38554 7972 38898
rect 7932 38548 7984 38554
rect 7932 38490 7984 38496
rect 8312 38350 8340 41398
rect 9600 40118 9628 42706
rect 11348 42702 11376 43046
rect 12452 42906 12480 43182
rect 12440 42900 12492 42906
rect 12440 42842 12492 42848
rect 12636 42702 12664 43590
rect 12716 43104 12768 43110
rect 12716 43046 12768 43052
rect 11336 42696 11388 42702
rect 11336 42638 11388 42644
rect 12624 42696 12676 42702
rect 12624 42638 12676 42644
rect 12728 42566 12756 43046
rect 12820 42702 12848 43590
rect 12992 43308 13044 43314
rect 12992 43250 13044 43256
rect 13004 42906 13032 43250
rect 12992 42900 13044 42906
rect 12992 42842 13044 42848
rect 12808 42696 12860 42702
rect 12808 42638 12860 42644
rect 12716 42560 12768 42566
rect 12716 42502 12768 42508
rect 12992 42560 13044 42566
rect 12992 42502 13044 42508
rect 13004 42226 13032 42502
rect 12992 42220 13044 42226
rect 12992 42162 13044 42168
rect 12624 42016 12676 42022
rect 12624 41958 12676 41964
rect 9588 40112 9640 40118
rect 9588 40054 9640 40060
rect 9312 39976 9364 39982
rect 9312 39918 9364 39924
rect 8484 39840 8536 39846
rect 8484 39782 8536 39788
rect 8496 39438 8524 39782
rect 8484 39432 8536 39438
rect 8484 39374 8536 39380
rect 8944 39432 8996 39438
rect 8944 39374 8996 39380
rect 8956 39030 8984 39374
rect 9324 39098 9352 39918
rect 9600 39438 9628 40054
rect 12636 40050 12664 41958
rect 11060 40044 11112 40050
rect 11060 39986 11112 39992
rect 12072 40044 12124 40050
rect 12072 39986 12124 39992
rect 12624 40044 12676 40050
rect 12624 39986 12676 39992
rect 11072 39642 11100 39986
rect 11060 39636 11112 39642
rect 11060 39578 11112 39584
rect 9588 39432 9640 39438
rect 9588 39374 9640 39380
rect 9312 39092 9364 39098
rect 9312 39034 9364 39040
rect 8944 39024 8996 39030
rect 8944 38966 8996 38972
rect 8300 38344 8352 38350
rect 8576 38344 8628 38350
rect 8352 38304 8524 38332
rect 8300 38286 8352 38292
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 8496 37806 8524 38304
rect 8576 38286 8628 38292
rect 8588 38010 8616 38286
rect 8576 38004 8628 38010
rect 8576 37946 8628 37952
rect 9324 37942 9352 39034
rect 9600 38962 9628 39374
rect 9680 39296 9732 39302
rect 9680 39238 9732 39244
rect 10324 39296 10376 39302
rect 10324 39238 10376 39244
rect 9588 38956 9640 38962
rect 9588 38898 9640 38904
rect 9692 38350 9720 39238
rect 9864 38956 9916 38962
rect 9864 38898 9916 38904
rect 9876 38554 9904 38898
rect 9864 38548 9916 38554
rect 9864 38490 9916 38496
rect 9680 38344 9732 38350
rect 9680 38286 9732 38292
rect 10336 38282 10364 39238
rect 10600 38752 10652 38758
rect 10600 38694 10652 38700
rect 10612 38350 10640 38694
rect 10600 38344 10652 38350
rect 10600 38286 10652 38292
rect 10324 38276 10376 38282
rect 10324 38218 10376 38224
rect 10140 38208 10192 38214
rect 10140 38150 10192 38156
rect 9312 37936 9364 37942
rect 9312 37878 9364 37884
rect 8484 37800 8536 37806
rect 8484 37742 8536 37748
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 8300 37460 8352 37466
rect 8300 37402 8352 37408
rect 8024 37188 8076 37194
rect 8024 37130 8076 37136
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 8036 36922 8064 37130
rect 8024 36916 8076 36922
rect 8024 36858 8076 36864
rect 8312 36650 8340 37402
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 8300 36644 8352 36650
rect 8300 36586 8352 36592
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 6920 35828 6972 35834
rect 6920 35770 6972 35776
rect 6368 35624 6420 35630
rect 6368 35566 6420 35572
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 6380 35290 6408 35566
rect 6368 35284 6420 35290
rect 6368 35226 6420 35232
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4620 34536 4672 34542
rect 4620 34478 4672 34484
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 33658 4660 34478
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4620 33652 4672 33658
rect 4620 33594 4672 33600
rect 3516 33516 3568 33522
rect 3516 33458 3568 33464
rect 2964 33448 3016 33454
rect 2964 33390 3016 33396
rect 848 32904 900 32910
rect 846 32872 848 32881
rect 900 32872 902 32881
rect 846 32807 902 32816
rect 848 32224 900 32230
rect 846 32192 848 32201
rect 900 32192 902 32201
rect 846 32127 902 32136
rect 848 31816 900 31822
rect 848 31758 900 31764
rect 860 31521 888 31758
rect 846 31512 902 31521
rect 846 31447 902 31456
rect 846 30832 902 30841
rect 846 30767 848 30776
rect 900 30767 902 30776
rect 848 30738 900 30744
rect 2976 30734 3004 33390
rect 3528 33114 3556 33458
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 6932 31346 6960 35770
rect 8312 35154 8340 36586
rect 8404 35766 8432 37198
rect 8496 36786 8524 37742
rect 9324 37330 9352 37878
rect 9680 37868 9732 37874
rect 9680 37810 9732 37816
rect 9692 37398 9720 37810
rect 9772 37664 9824 37670
rect 9772 37606 9824 37612
rect 9680 37392 9732 37398
rect 9680 37334 9732 37340
rect 9312 37324 9364 37330
rect 9312 37266 9364 37272
rect 9692 37262 9720 37334
rect 9220 37256 9272 37262
rect 9220 37198 9272 37204
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 8484 36780 8536 36786
rect 8484 36722 8536 36728
rect 9232 36242 9260 37198
rect 9312 37188 9364 37194
rect 9312 37130 9364 37136
rect 9324 36718 9352 37130
rect 9784 36786 9812 37606
rect 10152 37466 10180 38150
rect 10336 37942 10364 38218
rect 10612 38010 10640 38286
rect 10600 38004 10652 38010
rect 10600 37946 10652 37952
rect 10324 37936 10376 37942
rect 10324 37878 10376 37884
rect 10140 37460 10192 37466
rect 10140 37402 10192 37408
rect 10336 37330 10364 37878
rect 10508 37664 10560 37670
rect 10508 37606 10560 37612
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 10520 36854 10548 37606
rect 11072 37194 11100 39578
rect 12084 39506 12112 39986
rect 12072 39500 12124 39506
rect 12072 39442 12124 39448
rect 12440 39432 12492 39438
rect 12440 39374 12492 39380
rect 12256 39364 12308 39370
rect 12256 39306 12308 39312
rect 11152 37800 11204 37806
rect 11152 37742 11204 37748
rect 10968 37188 11020 37194
rect 10968 37130 11020 37136
rect 11060 37188 11112 37194
rect 11060 37130 11112 37136
rect 10980 36922 11008 37130
rect 11164 37126 11192 37742
rect 11152 37120 11204 37126
rect 11152 37062 11204 37068
rect 10968 36916 11020 36922
rect 10968 36858 11020 36864
rect 10508 36848 10560 36854
rect 10508 36790 10560 36796
rect 11796 36848 11848 36854
rect 11796 36790 11848 36796
rect 9772 36780 9824 36786
rect 9772 36722 9824 36728
rect 9312 36712 9364 36718
rect 9312 36654 9364 36660
rect 9680 36712 9732 36718
rect 9680 36654 9732 36660
rect 9220 36236 9272 36242
rect 9220 36178 9272 36184
rect 8944 36032 8996 36038
rect 8944 35974 8996 35980
rect 8392 35760 8444 35766
rect 8392 35702 8444 35708
rect 7012 35148 7064 35154
rect 7012 35090 7064 35096
rect 8300 35148 8352 35154
rect 8300 35090 8352 35096
rect 7024 34746 7052 35090
rect 8404 35018 8432 35702
rect 8956 35698 8984 35974
rect 9324 35834 9352 36654
rect 9496 36236 9548 36242
rect 9496 36178 9548 36184
rect 9312 35828 9364 35834
rect 9312 35770 9364 35776
rect 8944 35692 8996 35698
rect 8944 35634 8996 35640
rect 9508 35562 9536 36178
rect 9692 35766 9720 36654
rect 9680 35760 9732 35766
rect 9680 35702 9732 35708
rect 9496 35556 9548 35562
rect 9496 35498 9548 35504
rect 8392 35012 8444 35018
rect 8392 34954 8444 34960
rect 8852 34944 8904 34950
rect 8852 34886 8904 34892
rect 7012 34740 7064 34746
rect 7012 34682 7064 34688
rect 8864 34542 8892 34886
rect 9692 34678 9720 35702
rect 10692 35624 10744 35630
rect 10692 35566 10744 35572
rect 10704 34950 10732 35566
rect 11808 35290 11836 36790
rect 12268 36106 12296 39306
rect 12452 37942 12480 39374
rect 13188 39370 13216 43726
rect 13832 43450 13860 43726
rect 14660 43450 14688 43726
rect 13360 43444 13412 43450
rect 13360 43386 13412 43392
rect 13820 43444 13872 43450
rect 13820 43386 13872 43392
rect 14648 43444 14700 43450
rect 14648 43386 14700 43392
rect 13268 42696 13320 42702
rect 13268 42638 13320 42644
rect 13176 39364 13228 39370
rect 13176 39306 13228 39312
rect 13188 39098 13216 39306
rect 13176 39092 13228 39098
rect 13176 39034 13228 39040
rect 12532 38344 12584 38350
rect 12532 38286 12584 38292
rect 12440 37936 12492 37942
rect 12440 37878 12492 37884
rect 12440 37188 12492 37194
rect 12440 37130 12492 37136
rect 12452 36922 12480 37130
rect 12544 37126 12572 38286
rect 12624 37936 12676 37942
rect 12624 37878 12676 37884
rect 12532 37120 12584 37126
rect 12532 37062 12584 37068
rect 12440 36916 12492 36922
rect 12440 36858 12492 36864
rect 12544 36786 12572 37062
rect 12636 36854 12664 37878
rect 13280 37874 13308 42638
rect 13372 39438 13400 43386
rect 22836 43376 22888 43382
rect 22836 43318 22888 43324
rect 20168 43308 20220 43314
rect 20168 43250 20220 43256
rect 20180 41818 20208 43250
rect 21272 43104 21324 43110
rect 21272 43046 21324 43052
rect 21284 42770 21312 43046
rect 21272 42764 21324 42770
rect 21272 42706 21324 42712
rect 20812 42560 20864 42566
rect 20812 42502 20864 42508
rect 20168 41812 20220 41818
rect 20168 41754 20220 41760
rect 20824 41614 20852 42502
rect 17132 41608 17184 41614
rect 17132 41550 17184 41556
rect 20168 41608 20220 41614
rect 20168 41550 20220 41556
rect 20628 41608 20680 41614
rect 20628 41550 20680 41556
rect 20812 41608 20864 41614
rect 20812 41550 20864 41556
rect 16672 41540 16724 41546
rect 16672 41482 16724 41488
rect 16684 41274 16712 41482
rect 17040 41472 17092 41478
rect 17040 41414 17092 41420
rect 16672 41268 16724 41274
rect 16672 41210 16724 41216
rect 16580 41200 16632 41206
rect 16580 41142 16632 41148
rect 13452 39840 13504 39846
rect 13452 39782 13504 39788
rect 13360 39432 13412 39438
rect 13360 39374 13412 39380
rect 13372 38962 13400 39374
rect 13464 38962 13492 39782
rect 16212 39364 16264 39370
rect 16212 39306 16264 39312
rect 14556 39296 14608 39302
rect 14556 39238 14608 39244
rect 14568 38962 14596 39238
rect 16224 39098 16252 39306
rect 16212 39092 16264 39098
rect 16212 39034 16264 39040
rect 13360 38956 13412 38962
rect 13360 38898 13412 38904
rect 13452 38956 13504 38962
rect 13452 38898 13504 38904
rect 14556 38956 14608 38962
rect 14556 38898 14608 38904
rect 16028 38956 16080 38962
rect 16028 38898 16080 38904
rect 16212 38956 16264 38962
rect 16212 38898 16264 38904
rect 13464 38418 13492 38898
rect 14280 38888 14332 38894
rect 14280 38830 14332 38836
rect 14292 38554 14320 38830
rect 14280 38548 14332 38554
rect 14280 38490 14332 38496
rect 13452 38412 13504 38418
rect 13452 38354 13504 38360
rect 13268 37868 13320 37874
rect 13268 37810 13320 37816
rect 13464 37806 13492 38354
rect 13728 38344 13780 38350
rect 13728 38286 13780 38292
rect 13740 37874 13768 38286
rect 14292 38214 14320 38490
rect 14568 38350 14596 38898
rect 15384 38752 15436 38758
rect 15384 38694 15436 38700
rect 15396 38350 15424 38694
rect 16040 38486 16068 38898
rect 16028 38480 16080 38486
rect 16028 38422 16080 38428
rect 14556 38344 14608 38350
rect 14556 38286 14608 38292
rect 14648 38344 14700 38350
rect 14648 38286 14700 38292
rect 15384 38344 15436 38350
rect 15384 38286 15436 38292
rect 14280 38208 14332 38214
rect 14280 38150 14332 38156
rect 14292 37874 14320 38150
rect 14568 37942 14596 38286
rect 14556 37936 14608 37942
rect 14556 37878 14608 37884
rect 14660 37874 14688 38286
rect 16040 38010 16068 38422
rect 16224 38214 16252 38898
rect 16592 38758 16620 41142
rect 17052 41070 17080 41414
rect 17040 41064 17092 41070
rect 17040 41006 17092 41012
rect 17052 39506 17080 41006
rect 16764 39500 16816 39506
rect 16764 39442 16816 39448
rect 17040 39500 17092 39506
rect 17040 39442 17092 39448
rect 16580 38752 16632 38758
rect 16580 38694 16632 38700
rect 16672 38752 16724 38758
rect 16672 38694 16724 38700
rect 16684 38554 16712 38694
rect 16776 38554 16804 39442
rect 16856 39092 16908 39098
rect 16856 39034 16908 39040
rect 16868 38554 16896 39034
rect 17144 39030 17172 41550
rect 19616 41200 19668 41206
rect 19616 41142 19668 41148
rect 17592 41132 17644 41138
rect 17592 41074 17644 41080
rect 17604 40934 17632 41074
rect 17592 40928 17644 40934
rect 17592 40870 17644 40876
rect 17604 40526 17632 40870
rect 17592 40520 17644 40526
rect 17592 40462 17644 40468
rect 17604 39642 17632 40462
rect 17408 39636 17460 39642
rect 17408 39578 17460 39584
rect 17592 39636 17644 39642
rect 17592 39578 17644 39584
rect 18328 39636 18380 39642
rect 18328 39578 18380 39584
rect 17224 39296 17276 39302
rect 17224 39238 17276 39244
rect 17132 39024 17184 39030
rect 17132 38966 17184 38972
rect 16672 38548 16724 38554
rect 16672 38490 16724 38496
rect 16764 38548 16816 38554
rect 16764 38490 16816 38496
rect 16856 38548 16908 38554
rect 16856 38490 16908 38496
rect 17236 38418 17264 39238
rect 17420 38418 17448 39578
rect 17776 39364 17828 39370
rect 17776 39306 17828 39312
rect 17788 38758 17816 39306
rect 18340 38962 18368 39578
rect 18512 39296 18564 39302
rect 18512 39238 18564 39244
rect 19432 39296 19484 39302
rect 19432 39238 19484 39244
rect 18328 38956 18380 38962
rect 18328 38898 18380 38904
rect 18524 38944 18552 39238
rect 19444 39098 19472 39238
rect 19432 39092 19484 39098
rect 19432 39034 19484 39040
rect 19524 39024 19576 39030
rect 19524 38966 19576 38972
rect 18604 38956 18656 38962
rect 18524 38916 18604 38944
rect 18236 38820 18288 38826
rect 18236 38762 18288 38768
rect 17776 38752 17828 38758
rect 17776 38694 17828 38700
rect 18144 38752 18196 38758
rect 18144 38694 18196 38700
rect 17224 38412 17276 38418
rect 17224 38354 17276 38360
rect 17408 38412 17460 38418
rect 17408 38354 17460 38360
rect 16948 38344 17000 38350
rect 16948 38286 17000 38292
rect 17684 38344 17736 38350
rect 17684 38286 17736 38292
rect 16212 38208 16264 38214
rect 16212 38150 16264 38156
rect 16488 38208 16540 38214
rect 16488 38150 16540 38156
rect 16028 38004 16080 38010
rect 16028 37946 16080 37952
rect 13728 37868 13780 37874
rect 13728 37810 13780 37816
rect 14280 37868 14332 37874
rect 14280 37810 14332 37816
rect 14648 37868 14700 37874
rect 14648 37810 14700 37816
rect 12716 37800 12768 37806
rect 12716 37742 12768 37748
rect 13452 37800 13504 37806
rect 13452 37742 13504 37748
rect 12624 36848 12676 36854
rect 12624 36790 12676 36796
rect 12532 36780 12584 36786
rect 12532 36722 12584 36728
rect 12256 36100 12308 36106
rect 12256 36042 12308 36048
rect 12268 35894 12296 36042
rect 12728 35894 12756 37742
rect 14292 37126 14320 37810
rect 16500 37806 16528 38150
rect 16488 37800 16540 37806
rect 16488 37742 16540 37748
rect 16960 37670 16988 38286
rect 17696 38010 17724 38286
rect 17788 38010 17816 38694
rect 18156 38486 18184 38694
rect 18144 38480 18196 38486
rect 18144 38422 18196 38428
rect 18248 38350 18276 38762
rect 18236 38344 18288 38350
rect 18236 38286 18288 38292
rect 18328 38208 18380 38214
rect 18328 38150 18380 38156
rect 17684 38004 17736 38010
rect 17684 37946 17736 37952
rect 17776 38004 17828 38010
rect 17776 37946 17828 37952
rect 18340 37942 18368 38150
rect 18328 37936 18380 37942
rect 18328 37878 18380 37884
rect 16948 37664 17000 37670
rect 16948 37606 17000 37612
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 12176 35866 12296 35894
rect 12636 35866 12756 35894
rect 12072 35760 12124 35766
rect 12072 35702 12124 35708
rect 11888 35692 11940 35698
rect 11888 35634 11940 35640
rect 11900 35290 11928 35634
rect 11796 35284 11848 35290
rect 11796 35226 11848 35232
rect 11888 35284 11940 35290
rect 11888 35226 11940 35232
rect 12084 35086 12112 35702
rect 11152 35080 11204 35086
rect 11152 35022 11204 35028
rect 12072 35080 12124 35086
rect 12072 35022 12124 35028
rect 10692 34944 10744 34950
rect 10692 34886 10744 34892
rect 11164 34746 11192 35022
rect 12176 35018 12204 35866
rect 12164 35012 12216 35018
rect 12164 34954 12216 34960
rect 11152 34740 11204 34746
rect 11152 34682 11204 34688
rect 9680 34672 9732 34678
rect 9680 34614 9732 34620
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8864 33454 8892 34478
rect 8852 33448 8904 33454
rect 8852 33390 8904 33396
rect 8864 31822 8892 33390
rect 12532 33040 12584 33046
rect 12532 32982 12584 32988
rect 11888 32904 11940 32910
rect 11888 32846 11940 32852
rect 12440 32904 12492 32910
rect 12440 32846 12492 32852
rect 8852 31816 8904 31822
rect 8852 31758 8904 31764
rect 11704 31816 11756 31822
rect 11704 31758 11756 31764
rect 8668 31748 8720 31754
rect 8668 31690 8720 31696
rect 8680 31482 8708 31690
rect 8668 31476 8720 31482
rect 8668 31418 8720 31424
rect 8576 31408 8628 31414
rect 8576 31350 8628 31356
rect 6920 31340 6972 31346
rect 6920 31282 6972 31288
rect 5816 31272 5868 31278
rect 5816 31214 5868 31220
rect 6460 31272 6512 31278
rect 6460 31214 6512 31220
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 2964 30728 3016 30734
rect 2964 30670 3016 30676
rect 2976 29646 3004 30670
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5460 30258 5488 31078
rect 5448 30252 5500 30258
rect 5448 30194 5500 30200
rect 4712 30184 4764 30190
rect 4712 30126 4764 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4724 29646 4752 30126
rect 848 29640 900 29646
rect 848 29582 900 29588
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 4712 29640 4764 29646
rect 4712 29582 4764 29588
rect 860 29481 888 29582
rect 846 29472 902 29481
rect 846 29407 902 29416
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 5828 29306 5856 31214
rect 6368 31136 6420 31142
rect 6368 31078 6420 31084
rect 6380 29578 6408 31078
rect 6472 30938 6500 31214
rect 6460 30932 6512 30938
rect 6460 30874 6512 30880
rect 6932 30802 6960 31282
rect 6920 30796 6972 30802
rect 6920 30738 6972 30744
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 6736 30728 6788 30734
rect 6736 30670 6788 30676
rect 6932 30682 6960 30738
rect 6644 30592 6696 30598
rect 6644 30534 6696 30540
rect 6656 30326 6684 30534
rect 6644 30320 6696 30326
rect 6644 30262 6696 30268
rect 6748 29782 6776 30670
rect 6932 30654 7052 30682
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 6932 29866 6960 30534
rect 7024 30258 7052 30654
rect 7012 30252 7064 30258
rect 7012 30194 7064 30200
rect 7116 30054 7144 30738
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 7104 30048 7156 30054
rect 7104 29990 7156 29996
rect 7288 30048 7340 30054
rect 7288 29990 7340 29996
rect 6840 29850 6960 29866
rect 6828 29844 6960 29850
rect 6880 29838 6960 29844
rect 6828 29786 6880 29792
rect 6736 29776 6788 29782
rect 6736 29718 6788 29724
rect 6748 29578 6776 29718
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6736 29572 6788 29578
rect 6736 29514 6788 29520
rect 5816 29300 5868 29306
rect 5816 29242 5868 29248
rect 6932 29170 6960 29838
rect 7116 29646 7144 29990
rect 7104 29640 7156 29646
rect 7104 29582 7156 29588
rect 7300 29170 7328 29990
rect 7392 29170 7420 30194
rect 7748 30116 7800 30122
rect 7748 30058 7800 30064
rect 7760 29850 7788 30058
rect 7748 29844 7800 29850
rect 7748 29786 7800 29792
rect 7656 29572 7708 29578
rect 7656 29514 7708 29520
rect 7668 29306 7696 29514
rect 7656 29300 7708 29306
rect 7656 29242 7708 29248
rect 8588 29170 8616 31350
rect 8864 30326 8892 31758
rect 10324 31680 10376 31686
rect 10324 31622 10376 31628
rect 9220 31272 9272 31278
rect 9220 31214 9272 31220
rect 9232 30666 9260 31214
rect 9588 30728 9640 30734
rect 9588 30670 9640 30676
rect 9220 30660 9272 30666
rect 9220 30602 9272 30608
rect 8944 30592 8996 30598
rect 8944 30534 8996 30540
rect 8852 30320 8904 30326
rect 8852 30262 8904 30268
rect 8864 29646 8892 30262
rect 8956 29714 8984 30534
rect 9232 30054 9260 30602
rect 9600 30326 9628 30670
rect 9588 30320 9640 30326
rect 9588 30262 9640 30268
rect 9220 30048 9272 30054
rect 9220 29990 9272 29996
rect 8944 29708 8996 29714
rect 8944 29650 8996 29656
rect 8852 29640 8904 29646
rect 8852 29582 8904 29588
rect 8668 29504 8720 29510
rect 8668 29446 8720 29452
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 7288 29164 7340 29170
rect 7288 29106 7340 29112
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 8576 29164 8628 29170
rect 8576 29106 8628 29112
rect 8680 29102 8708 29446
rect 8864 29170 8892 29582
rect 9232 29238 9260 29990
rect 9496 29640 9548 29646
rect 9496 29582 9548 29588
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9220 29232 9272 29238
rect 9220 29174 9272 29180
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 8668 29096 8720 29102
rect 8668 29038 8720 29044
rect 848 29028 900 29034
rect 848 28970 900 28976
rect 860 28801 888 28970
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 846 28792 902 28801
rect 4214 28795 4522 28804
rect 846 28727 902 28736
rect 9416 28558 9444 29446
rect 9508 28558 9536 29582
rect 10336 29578 10364 31622
rect 11716 31346 11744 31758
rect 11900 31346 11928 32846
rect 12452 32230 12480 32846
rect 12544 32366 12572 32982
rect 12636 32910 12664 35866
rect 18340 35018 18368 37878
rect 18328 35012 18380 35018
rect 18328 34954 18380 34960
rect 18340 34678 18368 34954
rect 18328 34672 18380 34678
rect 18328 34614 18380 34620
rect 18524 34610 18552 38916
rect 18604 38898 18656 38904
rect 18880 38888 18932 38894
rect 18880 38830 18932 38836
rect 18696 38752 18748 38758
rect 18696 38694 18748 38700
rect 18708 38418 18736 38694
rect 18696 38412 18748 38418
rect 18696 38354 18748 38360
rect 18892 38282 18920 38830
rect 19340 38752 19392 38758
rect 19340 38694 19392 38700
rect 18880 38276 18932 38282
rect 18880 38218 18932 38224
rect 19352 36786 19380 38694
rect 19536 38554 19564 38966
rect 19524 38548 19576 38554
rect 19524 38490 19576 38496
rect 19628 38282 19656 41142
rect 20180 41138 20208 41550
rect 20536 41540 20588 41546
rect 20536 41482 20588 41488
rect 20168 41132 20220 41138
rect 20168 41074 20220 41080
rect 20548 40730 20576 41482
rect 20536 40724 20588 40730
rect 20536 40666 20588 40672
rect 20640 40662 20668 41550
rect 21088 41472 21140 41478
rect 21088 41414 21140 41420
rect 21100 40730 21128 41414
rect 21180 40996 21232 41002
rect 21180 40938 21232 40944
rect 21088 40724 21140 40730
rect 21088 40666 21140 40672
rect 21192 40662 21220 40938
rect 20628 40656 20680 40662
rect 20628 40598 20680 40604
rect 21180 40656 21232 40662
rect 21180 40598 21232 40604
rect 21088 40588 21140 40594
rect 21088 40530 21140 40536
rect 20996 40520 21048 40526
rect 20996 40462 21048 40468
rect 21008 40186 21036 40462
rect 20996 40180 21048 40186
rect 20996 40122 21048 40128
rect 19892 40044 19944 40050
rect 19892 39986 19944 39992
rect 20076 40044 20128 40050
rect 20076 39986 20128 39992
rect 20812 40044 20864 40050
rect 20812 39986 20864 39992
rect 20996 40044 21048 40050
rect 20996 39986 21048 39992
rect 19800 39840 19852 39846
rect 19800 39782 19852 39788
rect 19812 39438 19840 39782
rect 19904 39438 19932 39986
rect 20088 39438 20116 39986
rect 20168 39908 20220 39914
rect 20168 39850 20220 39856
rect 20180 39642 20208 39850
rect 20444 39840 20496 39846
rect 20444 39782 20496 39788
rect 20628 39840 20680 39846
rect 20628 39782 20680 39788
rect 20168 39636 20220 39642
rect 20168 39578 20220 39584
rect 20456 39506 20484 39782
rect 20444 39500 20496 39506
rect 20444 39442 20496 39448
rect 19800 39432 19852 39438
rect 19800 39374 19852 39380
rect 19892 39432 19944 39438
rect 19892 39374 19944 39380
rect 20076 39432 20128 39438
rect 20076 39374 20128 39380
rect 19904 38962 19932 39374
rect 19892 38956 19944 38962
rect 19892 38898 19944 38904
rect 20088 38554 20116 39374
rect 20260 38956 20312 38962
rect 20260 38898 20312 38904
rect 20076 38548 20128 38554
rect 20076 38490 20128 38496
rect 19616 38276 19668 38282
rect 19616 38218 19668 38224
rect 19628 38010 19656 38218
rect 20272 38214 20300 38898
rect 20444 38820 20496 38826
rect 20444 38762 20496 38768
rect 20456 38350 20484 38762
rect 20536 38752 20588 38758
rect 20536 38694 20588 38700
rect 20548 38486 20576 38694
rect 20536 38480 20588 38486
rect 20536 38422 20588 38428
rect 20640 38418 20668 39782
rect 20824 38826 20852 39986
rect 21008 39642 21036 39986
rect 21100 39642 21128 40530
rect 20996 39636 21048 39642
rect 20996 39578 21048 39584
rect 21088 39636 21140 39642
rect 21088 39578 21140 39584
rect 21192 38894 21220 40598
rect 21284 39914 21312 42706
rect 22848 41614 22876 43318
rect 22836 41608 22888 41614
rect 22836 41550 22888 41556
rect 21364 40044 21416 40050
rect 21364 39986 21416 39992
rect 21272 39908 21324 39914
rect 21272 39850 21324 39856
rect 21376 39846 21404 39986
rect 21640 39908 21692 39914
rect 21640 39850 21692 39856
rect 21364 39840 21416 39846
rect 21364 39782 21416 39788
rect 21272 39636 21324 39642
rect 21376 39624 21404 39782
rect 21324 39596 21404 39624
rect 21272 39578 21324 39584
rect 21284 39506 21312 39578
rect 21272 39500 21324 39506
rect 21272 39442 21324 39448
rect 21652 39438 21680 39850
rect 21364 39432 21416 39438
rect 21364 39374 21416 39380
rect 21640 39432 21692 39438
rect 21640 39374 21692 39380
rect 21180 38888 21232 38894
rect 21180 38830 21232 38836
rect 20812 38820 20864 38826
rect 20812 38762 20864 38768
rect 20628 38412 20680 38418
rect 20628 38354 20680 38360
rect 20444 38344 20496 38350
rect 20444 38286 20496 38292
rect 20260 38208 20312 38214
rect 20260 38150 20312 38156
rect 19616 38004 19668 38010
rect 19616 37946 19668 37952
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 19892 36100 19944 36106
rect 19892 36042 19944 36048
rect 18604 35760 18656 35766
rect 18604 35702 18656 35708
rect 18616 34610 18644 35702
rect 18880 35692 18932 35698
rect 18880 35634 18932 35640
rect 18892 35222 18920 35634
rect 18880 35216 18932 35222
rect 18880 35158 18932 35164
rect 18892 34610 18920 35158
rect 19524 35148 19576 35154
rect 19524 35090 19576 35096
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 19340 34944 19392 34950
rect 19340 34886 19392 34892
rect 16212 34604 16264 34610
rect 16212 34546 16264 34552
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 18604 34604 18656 34610
rect 18604 34546 18656 34552
rect 18880 34604 18932 34610
rect 18880 34546 18932 34552
rect 15016 34400 15068 34406
rect 15016 34342 15068 34348
rect 15028 33998 15056 34342
rect 16224 34202 16252 34546
rect 17776 34536 17828 34542
rect 17776 34478 17828 34484
rect 17788 34202 17816 34478
rect 16212 34196 16264 34202
rect 16212 34138 16264 34144
rect 17776 34196 17828 34202
rect 17776 34138 17828 34144
rect 17500 34060 17552 34066
rect 17500 34002 17552 34008
rect 15016 33992 15068 33998
rect 15016 33934 15068 33940
rect 16672 33992 16724 33998
rect 16672 33934 16724 33940
rect 15028 33522 15056 33934
rect 15108 33924 15160 33930
rect 15108 33866 15160 33872
rect 15120 33522 15148 33866
rect 15936 33856 15988 33862
rect 15936 33798 15988 33804
rect 15476 33584 15528 33590
rect 15476 33526 15528 33532
rect 13268 33516 13320 33522
rect 13268 33458 13320 33464
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 15108 33516 15160 33522
rect 15108 33458 15160 33464
rect 13280 33114 13308 33458
rect 13912 33380 13964 33386
rect 13912 33322 13964 33328
rect 13268 33108 13320 33114
rect 13268 33050 13320 33056
rect 13636 33108 13688 33114
rect 13636 33050 13688 33056
rect 12900 32972 12952 32978
rect 12900 32914 12952 32920
rect 12624 32904 12676 32910
rect 12624 32846 12676 32852
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 11980 32224 12032 32230
rect 11980 32166 12032 32172
rect 12440 32224 12492 32230
rect 12440 32166 12492 32172
rect 11992 31346 12020 32166
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11980 31340 12032 31346
rect 11980 31282 12032 31288
rect 12440 31340 12492 31346
rect 12440 31282 12492 31288
rect 11520 31136 11572 31142
rect 11520 31078 11572 31084
rect 11532 30734 11560 31078
rect 11520 30728 11572 30734
rect 11520 30670 11572 30676
rect 11900 30394 11928 31282
rect 12452 30410 12480 31282
rect 12544 30938 12572 32302
rect 12636 31346 12664 32846
rect 12912 32570 12940 32914
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 12808 32428 12860 32434
rect 12808 32370 12860 32376
rect 12716 31884 12768 31890
rect 12716 31826 12768 31832
rect 12728 31657 12756 31826
rect 12714 31648 12770 31657
rect 12714 31583 12770 31592
rect 12820 31482 12848 32370
rect 12912 31822 12940 32506
rect 13648 32434 13676 33050
rect 13820 32768 13872 32774
rect 13820 32710 13872 32716
rect 13832 32502 13860 32710
rect 13820 32496 13872 32502
rect 13820 32438 13872 32444
rect 13924 32434 13952 33322
rect 14004 33312 14056 33318
rect 14004 33254 14056 33260
rect 14016 32910 14044 33254
rect 15120 33114 15148 33458
rect 15292 33448 15344 33454
rect 15292 33390 15344 33396
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 14096 33040 14148 33046
rect 14096 32982 14148 32988
rect 14004 32904 14056 32910
rect 14004 32846 14056 32852
rect 14108 32434 14136 32982
rect 15304 32910 15332 33390
rect 15384 33380 15436 33386
rect 15384 33322 15436 33328
rect 15396 32910 15424 33322
rect 15488 32910 15516 33526
rect 15948 33386 15976 33798
rect 16684 33658 16712 33934
rect 16672 33652 16724 33658
rect 16672 33594 16724 33600
rect 17512 33522 17540 34002
rect 17592 33652 17644 33658
rect 17592 33594 17644 33600
rect 17500 33516 17552 33522
rect 17500 33458 17552 33464
rect 17224 33448 17276 33454
rect 17224 33390 17276 33396
rect 15936 33380 15988 33386
rect 15936 33322 15988 33328
rect 17236 32978 17264 33390
rect 16580 32972 16632 32978
rect 16580 32914 16632 32920
rect 17224 32972 17276 32978
rect 17224 32914 17276 32920
rect 15292 32904 15344 32910
rect 15292 32846 15344 32852
rect 15384 32904 15436 32910
rect 15384 32846 15436 32852
rect 15476 32904 15528 32910
rect 15476 32846 15528 32852
rect 14188 32836 14240 32842
rect 14188 32778 14240 32784
rect 14200 32434 14228 32778
rect 15304 32570 15332 32846
rect 15568 32768 15620 32774
rect 15568 32710 15620 32716
rect 15292 32564 15344 32570
rect 15292 32506 15344 32512
rect 13636 32428 13688 32434
rect 13636 32370 13688 32376
rect 13912 32428 13964 32434
rect 13912 32370 13964 32376
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 14188 32428 14240 32434
rect 14188 32370 14240 32376
rect 13084 32360 13136 32366
rect 13084 32302 13136 32308
rect 13176 32360 13228 32366
rect 13648 32314 13676 32370
rect 13176 32302 13228 32308
rect 12992 32292 13044 32298
rect 12992 32234 13044 32240
rect 13004 32026 13032 32234
rect 13096 32026 13124 32302
rect 12992 32020 13044 32026
rect 12992 31962 13044 31968
rect 13084 32020 13136 32026
rect 13084 31962 13136 31968
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 12808 31476 12860 31482
rect 12808 31418 12860 31424
rect 13096 31414 13124 31962
rect 12716 31408 12768 31414
rect 12716 31350 12768 31356
rect 13084 31408 13136 31414
rect 13084 31350 13136 31356
rect 12624 31340 12676 31346
rect 12624 31282 12676 31288
rect 12624 31204 12676 31210
rect 12624 31146 12676 31152
rect 12532 30932 12584 30938
rect 12532 30874 12584 30880
rect 12636 30598 12664 31146
rect 12728 30734 12756 31350
rect 13188 31346 13216 32302
rect 13556 32286 13676 32314
rect 13360 31884 13412 31890
rect 13360 31826 13412 31832
rect 13268 31680 13320 31686
rect 13268 31622 13320 31628
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 13176 31340 13228 31346
rect 13176 31282 13228 31288
rect 12808 31204 12860 31210
rect 12808 31146 12860 31152
rect 12716 30728 12768 30734
rect 12716 30670 12768 30676
rect 12624 30592 12676 30598
rect 12624 30534 12676 30540
rect 11888 30388 11940 30394
rect 11888 30330 11940 30336
rect 12360 30382 12480 30410
rect 10692 30184 10744 30190
rect 10692 30126 10744 30132
rect 10600 29708 10652 29714
rect 10600 29650 10652 29656
rect 10416 29640 10468 29646
rect 10416 29582 10468 29588
rect 10324 29572 10376 29578
rect 10324 29514 10376 29520
rect 9680 29504 9732 29510
rect 9680 29446 9732 29452
rect 9692 29306 9720 29446
rect 9680 29300 9732 29306
rect 9680 29242 9732 29248
rect 10336 28966 10364 29514
rect 10428 29306 10456 29582
rect 10416 29300 10468 29306
rect 10416 29242 10468 29248
rect 10612 29170 10640 29650
rect 10704 29510 10732 30126
rect 11336 30048 11388 30054
rect 11336 29990 11388 29996
rect 11348 29850 11376 29990
rect 11336 29844 11388 29850
rect 11336 29786 11388 29792
rect 12360 29646 12388 30382
rect 12624 30184 12676 30190
rect 12624 30126 12676 30132
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10324 28960 10376 28966
rect 10324 28902 10376 28908
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 8944 28416 8996 28422
rect 8944 28358 8996 28364
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 8956 27062 8984 28358
rect 8944 27056 8996 27062
rect 8944 26998 8996 27004
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 8956 26450 8984 26862
rect 8944 26444 8996 26450
rect 8944 26386 8996 26392
rect 8956 26234 8984 26386
rect 8772 26206 8984 26234
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 8772 25362 8800 26206
rect 9508 26042 9536 28494
rect 10704 28422 10732 29446
rect 10784 28960 10836 28966
rect 10784 28902 10836 28908
rect 10796 28490 10824 28902
rect 10784 28484 10836 28490
rect 10784 28426 10836 28432
rect 10692 28416 10744 28422
rect 10692 28358 10744 28364
rect 12636 26926 12664 30126
rect 12624 26920 12676 26926
rect 12624 26862 12676 26868
rect 10324 26784 10376 26790
rect 10324 26726 10376 26732
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 8760 25356 8812 25362
rect 8760 25298 8812 25304
rect 7012 25288 7064 25294
rect 7012 25230 7064 25236
rect 6368 25152 6420 25158
rect 6368 25094 6420 25100
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 848 24812 900 24818
rect 848 24754 900 24760
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 860 24721 888 24754
rect 2504 24744 2556 24750
rect 846 24712 902 24721
rect 2504 24686 2556 24692
rect 846 24647 902 24656
rect 2516 24206 2544 24686
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 2504 24200 2556 24206
rect 2504 24142 2556 24148
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4724 23186 4752 24754
rect 4816 24410 4844 24754
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 6092 24608 6144 24614
rect 6092 24550 6144 24556
rect 5460 24410 5488 24550
rect 4804 24404 4856 24410
rect 4804 24346 4856 24352
rect 5448 24404 5500 24410
rect 5448 24346 5500 24352
rect 5460 24274 5488 24346
rect 6104 24274 6132 24550
rect 6380 24342 6408 25094
rect 7024 24614 7052 25230
rect 7840 25220 7892 25226
rect 7840 25162 7892 25168
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7012 24608 7064 24614
rect 7012 24550 7064 24556
rect 6736 24404 6788 24410
rect 6736 24346 6788 24352
rect 6368 24336 6420 24342
rect 6368 24278 6420 24284
rect 5448 24268 5500 24274
rect 5448 24210 5500 24216
rect 6092 24268 6144 24274
rect 6092 24210 6144 24216
rect 6380 24206 6408 24278
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5920 23730 5948 24142
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 6012 23730 6040 24006
rect 6380 23866 6408 24142
rect 6368 23860 6420 23866
rect 6368 23802 6420 23808
rect 6748 23730 6776 24346
rect 7024 24138 7052 24550
rect 7012 24132 7064 24138
rect 7012 24074 7064 24080
rect 7288 24132 7340 24138
rect 7288 24074 7340 24080
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7208 23730 7236 24006
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 6000 23724 6052 23730
rect 6000 23666 6052 23672
rect 6736 23724 6788 23730
rect 6736 23666 6788 23672
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 6368 23656 6420 23662
rect 6368 23598 6420 23604
rect 6828 23656 6880 23662
rect 6828 23598 6880 23604
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 5368 19922 5396 23054
rect 5736 23050 5764 23462
rect 5724 23044 5776 23050
rect 5724 22986 5776 22992
rect 6380 22778 6408 23598
rect 6840 23118 6868 23598
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 7116 23118 7144 23462
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 6736 22976 6788 22982
rect 6736 22918 6788 22924
rect 6748 22778 6776 22918
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6840 22710 6868 23054
rect 7012 23044 7064 23050
rect 7012 22986 7064 22992
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6828 22704 6880 22710
rect 6828 22646 6880 22652
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6748 21962 6776 22578
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6840 22166 6868 22510
rect 6828 22160 6880 22166
rect 6828 22102 6880 22108
rect 6736 21956 6788 21962
rect 6736 21898 6788 21904
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 6380 20466 6408 21830
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5368 19446 5396 19858
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 5368 18834 5396 19382
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5644 18766 5672 20198
rect 6748 19854 6776 21898
rect 6840 20058 6868 22102
rect 6932 22098 6960 22714
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 7024 21146 7052 22986
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 7116 22166 7144 22918
rect 7300 22642 7328 24074
rect 7484 23866 7512 24754
rect 7852 24410 7880 25162
rect 8116 25152 8168 25158
rect 8116 25094 8168 25100
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 8128 24206 8156 25094
rect 8404 24750 8432 25298
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7472 23860 7524 23866
rect 7472 23802 7524 23808
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7484 22642 7512 22918
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7104 22160 7156 22166
rect 7104 22102 7156 22108
rect 7760 22030 7788 24006
rect 8312 23730 8340 24210
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 8116 23044 8168 23050
rect 8116 22986 8168 22992
rect 8128 22778 8156 22986
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8312 22642 8340 23666
rect 8404 23118 8432 24686
rect 9416 24274 9444 25842
rect 9508 24886 9536 25978
rect 10336 25906 10364 26726
rect 12636 26382 12664 26862
rect 12624 26376 12676 26382
rect 12544 26324 12624 26330
rect 12544 26318 12676 26324
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 12544 26302 12664 26318
rect 12268 26042 12296 26250
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 12360 25922 12388 26182
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 12268 25894 12388 25922
rect 12440 25900 12492 25906
rect 9496 24880 9548 24886
rect 9496 24822 9548 24828
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9784 23118 9812 23666
rect 9876 23662 9904 25842
rect 12268 25838 12296 25894
rect 12440 25842 12492 25848
rect 12256 25832 12308 25838
rect 12256 25774 12308 25780
rect 12348 25832 12400 25838
rect 12348 25774 12400 25780
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12176 25362 12204 25638
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 12268 25294 12296 25774
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 10140 24608 10192 24614
rect 10140 24550 10192 24556
rect 10152 23798 10180 24550
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 9864 23656 9916 23662
rect 9916 23616 9996 23644
rect 9864 23598 9916 23604
rect 9968 23186 9996 23616
rect 9956 23180 10008 23186
rect 9956 23122 10008 23128
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 8668 23044 8720 23050
rect 8668 22986 8720 22992
rect 8680 22710 8708 22986
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 8772 22710 8800 22918
rect 8668 22704 8720 22710
rect 8668 22646 8720 22652
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8300 22636 8352 22642
rect 8220 22596 8300 22624
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6196 19514 6224 19790
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6380 19514 6408 19722
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6932 19310 6960 19654
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7024 18970 7052 20878
rect 7208 19310 7236 21082
rect 8220 20398 8248 22596
rect 8300 22578 8352 22584
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 7392 19514 7420 20334
rect 8312 20262 8340 20810
rect 8956 20262 8984 23054
rect 9784 22642 9812 23054
rect 9968 22642 9996 23122
rect 10152 23050 10180 23734
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 10428 23322 10456 23666
rect 11428 23588 11480 23594
rect 11428 23530 11480 23536
rect 11244 23520 11296 23526
rect 11244 23462 11296 23468
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 10140 23044 10192 23050
rect 10140 22986 10192 22992
rect 10152 22642 10180 22986
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 10140 22636 10192 22642
rect 10428 22624 10456 23258
rect 11256 23118 11284 23462
rect 11440 23118 11468 23530
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 10612 22778 10640 23054
rect 11704 23044 11756 23050
rect 11704 22986 11756 22992
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 10508 22636 10560 22642
rect 10428 22596 10508 22624
rect 10140 22578 10192 22584
rect 10508 22578 10560 22584
rect 11716 22574 11744 22986
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 11808 22098 11836 22918
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 12268 21962 12296 25230
rect 12360 25158 12388 25774
rect 12452 25294 12480 25842
rect 12544 25294 12572 26302
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12636 25702 12664 25842
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12452 24342 12480 25230
rect 12544 24954 12572 25230
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 12440 24336 12492 24342
rect 12440 24278 12492 24284
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12360 22234 12388 22918
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 12360 21962 12388 22170
rect 12820 22094 12848 31146
rect 12912 30734 12940 31282
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 12912 27130 12940 30670
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 13004 26246 13032 26930
rect 13176 26852 13228 26858
rect 13176 26794 13228 26800
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 12992 26240 13044 26246
rect 12992 26182 13044 26188
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 12912 25362 12940 25842
rect 13004 25430 13032 25842
rect 13096 25838 13124 26726
rect 13188 26042 13216 26794
rect 13176 26036 13228 26042
rect 13176 25978 13228 25984
rect 13084 25832 13136 25838
rect 13084 25774 13136 25780
rect 12992 25424 13044 25430
rect 12992 25366 13044 25372
rect 13176 25424 13228 25430
rect 13176 25366 13228 25372
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 12728 22066 12848 22094
rect 12912 22094 12940 25298
rect 12912 22066 13124 22094
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12452 21622 12480 21966
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 9496 20528 9548 20534
rect 9496 20470 9548 20476
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 8956 19854 8984 20198
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 7380 19508 7432 19514
rect 7380 19450 7432 19456
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 8772 18290 8800 19110
rect 8864 18290 8892 19314
rect 8956 18834 8984 19790
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 9048 18426 9076 18634
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5552 16250 5580 16526
rect 7668 16454 7696 16526
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5828 16114 5856 16390
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 860 15881 888 16050
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3240 15904 3292 15910
rect 846 15872 902 15881
rect 3240 15846 3292 15852
rect 846 15807 902 15816
rect 3252 15502 3280 15846
rect 3436 15706 3464 15982
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 6012 15502 6040 16050
rect 6288 15570 6316 16390
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 7300 15502 7328 15846
rect 7668 15706 7696 16390
rect 8312 16250 8340 16526
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 8036 15366 8064 15574
rect 8312 15434 8340 16050
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8496 15570 8524 15914
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 7576 14618 7604 14962
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7852 14414 7880 15302
rect 8312 14414 8340 15370
rect 8496 15162 8524 15506
rect 8588 15502 8616 16186
rect 9508 16182 9536 20470
rect 12176 20398 12204 21286
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12452 20330 12480 20878
rect 12544 20398 12572 21966
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12544 19854 12572 20198
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9784 18086 9812 19246
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9876 17542 9904 18226
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9876 16590 9904 17478
rect 10244 17270 10272 17614
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9968 16726 9996 16934
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9968 16250 9996 16526
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 9048 15434 9076 15846
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8496 14482 8524 15098
rect 9048 14958 9076 15370
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 940 10056 992 10062
rect 940 9998 992 10004
rect 952 9625 980 9998
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 938 9616 994 9625
rect 938 9551 994 9560
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5828 9042 5856 9522
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5644 8634 5672 8842
rect 7300 8634 7328 9522
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7576 8498 7604 8774
rect 7852 8566 7880 14350
rect 9048 11694 9076 14894
rect 9692 14618 9720 14962
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 10244 14414 10272 17206
rect 10336 16114 10364 18566
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10520 16574 10548 18022
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10796 16726 10824 17614
rect 11348 17202 11376 18158
rect 11520 17264 11572 17270
rect 11520 17206 11572 17212
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10520 16546 10640 16574
rect 10612 16114 10640 16546
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10336 14822 10364 16050
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10520 15094 10548 15302
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10612 14958 10640 16050
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10704 15162 10732 15982
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10796 15026 10824 16662
rect 11164 16658 11192 16934
rect 11256 16794 11284 17138
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11072 15706 11100 16458
rect 11164 16250 11192 16458
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11348 15502 11376 17138
rect 11532 16658 11560 17206
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 16794 12204 16934
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11532 15502 11560 16390
rect 11624 15706 11652 16662
rect 12176 16182 12204 16730
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 10980 15162 11008 15438
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 9784 12238 9812 14350
rect 12084 13394 12112 15982
rect 12544 15706 12572 16526
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12544 15026 12572 15642
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11830 9628 12038
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9048 11150 9076 11630
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9232 10810 9260 11018
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8772 9450 8800 10542
rect 9324 9654 9352 11018
rect 9784 10742 9812 12174
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5460 2650 5488 8434
rect 9324 8430 9352 9590
rect 9784 9586 9812 10678
rect 10152 10266 10180 10678
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10428 9722 10456 9998
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9178 9444 9454
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9784 8634 9812 9522
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9876 8566 9904 9318
rect 9968 8974 9996 9590
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10152 9110 10180 9522
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9324 7886 9352 8366
rect 9968 8090 9996 8910
rect 10428 8906 10456 9658
rect 10520 9058 10548 11494
rect 11348 10674 11376 11494
rect 11532 10674 11560 12378
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 11354 11744 12174
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11716 10810 11744 11290
rect 12084 11218 12112 13330
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12636 12442 12664 13194
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10612 9178 10640 9930
rect 10704 9722 10732 9998
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10796 9586 10824 10066
rect 10980 9994 11008 10406
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 11072 9926 11100 10202
rect 11532 10130 11560 10610
rect 11900 10266 11928 10610
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 12084 10062 12112 11154
rect 12728 10742 12756 22066
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13004 21894 13032 21966
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 13004 21418 13032 21830
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12912 20466 12940 20878
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13004 20466 13032 20742
rect 13096 20466 13124 22066
rect 13188 20942 13216 25366
rect 13280 25294 13308 31622
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13280 23322 13308 25230
rect 13372 24818 13400 31826
rect 13556 31754 13584 32286
rect 13820 32224 13872 32230
rect 13820 32166 13872 32172
rect 14004 32224 14056 32230
rect 14004 32166 14056 32172
rect 13832 31754 13860 32166
rect 14016 31890 14044 32166
rect 14200 31958 14228 32370
rect 14188 31952 14240 31958
rect 14188 31894 14240 31900
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 13544 31748 13596 31754
rect 13544 31690 13596 31696
rect 13820 31748 13872 31754
rect 13820 31690 13872 31696
rect 13556 31657 13584 31690
rect 13542 31648 13598 31657
rect 13542 31583 13598 31592
rect 13556 30190 13584 31583
rect 13832 30598 13860 31690
rect 15580 30734 15608 32710
rect 16592 31822 16620 32914
rect 16304 31816 16356 31822
rect 16304 31758 16356 31764
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 15660 30796 15712 30802
rect 15660 30738 15712 30744
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 13820 30592 13872 30598
rect 13820 30534 13872 30540
rect 15108 30592 15160 30598
rect 15108 30534 15160 30540
rect 13636 30388 13688 30394
rect 13636 30330 13688 30336
rect 13544 30184 13596 30190
rect 13544 30126 13596 30132
rect 13648 27470 13676 30330
rect 15120 29170 15148 30534
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15304 29510 15332 30194
rect 15672 30190 15700 30738
rect 15936 30592 15988 30598
rect 15936 30534 15988 30540
rect 15948 30326 15976 30534
rect 15936 30320 15988 30326
rect 15936 30262 15988 30268
rect 16316 30258 16344 31758
rect 16304 30252 16356 30258
rect 16304 30194 16356 30200
rect 16396 30252 16448 30258
rect 16396 30194 16448 30200
rect 15660 30184 15712 30190
rect 16408 30138 16436 30194
rect 15660 30126 15712 30132
rect 16316 30110 16436 30138
rect 16212 30048 16264 30054
rect 16212 29990 16264 29996
rect 16224 29646 16252 29990
rect 16212 29640 16264 29646
rect 16212 29582 16264 29588
rect 16316 29510 16344 30110
rect 15292 29504 15344 29510
rect 15292 29446 15344 29452
rect 16304 29504 16356 29510
rect 16304 29446 16356 29452
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 16316 28490 16344 29446
rect 17500 29028 17552 29034
rect 17500 28970 17552 28976
rect 16304 28484 16356 28490
rect 16304 28426 16356 28432
rect 13452 27464 13504 27470
rect 13452 27406 13504 27412
rect 13636 27464 13688 27470
rect 13688 27424 13768 27452
rect 13636 27406 13688 27412
rect 13464 26042 13492 27406
rect 13740 26926 13768 27424
rect 16316 27402 16344 28426
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 16764 27600 16816 27606
rect 16764 27542 16816 27548
rect 16304 27396 16356 27402
rect 16304 27338 16356 27344
rect 14004 27328 14056 27334
rect 14004 27270 14056 27276
rect 14016 26994 14044 27270
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 13636 26920 13688 26926
rect 13636 26862 13688 26868
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13648 26586 13676 26862
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13452 26036 13504 26042
rect 13452 25978 13504 25984
rect 13740 25838 13768 26862
rect 13728 25832 13780 25838
rect 13648 25780 13728 25786
rect 13648 25774 13780 25780
rect 13648 25758 13768 25774
rect 13648 25702 13676 25758
rect 13636 25696 13688 25702
rect 13636 25638 13688 25644
rect 13728 25696 13780 25702
rect 13728 25638 13780 25644
rect 13648 25430 13676 25638
rect 13740 25498 13768 25638
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13636 25424 13688 25430
rect 13636 25366 13688 25372
rect 13832 25362 13860 26930
rect 14200 26586 14228 26930
rect 14464 26784 14516 26790
rect 14464 26726 14516 26732
rect 14188 26580 14240 26586
rect 14188 26522 14240 26528
rect 13912 26512 13964 26518
rect 13912 26454 13964 26460
rect 13820 25356 13872 25362
rect 13820 25298 13872 25304
rect 13924 25226 13952 26454
rect 14200 26382 14228 26522
rect 14476 26382 14504 26726
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 14372 26376 14424 26382
rect 14372 26318 14424 26324
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 13912 25220 13964 25226
rect 13912 25162 13964 25168
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 13372 23254 13400 24754
rect 13556 24274 13584 24890
rect 13924 24818 13952 25162
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13636 24676 13688 24682
rect 13636 24618 13688 24624
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 13648 24206 13676 24618
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13648 23730 13676 24142
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13360 23248 13412 23254
rect 13360 23190 13412 23196
rect 13820 21956 13872 21962
rect 13820 21898 13872 21904
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 13188 20058 13216 20878
rect 13832 20534 13860 21898
rect 14384 20534 14412 26318
rect 16316 25906 16344 27338
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 16304 25900 16356 25906
rect 16304 25842 16356 25848
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15304 22778 15332 23666
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14660 21962 14688 22578
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 14372 20528 14424 20534
rect 14372 20470 14424 20476
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13280 19938 13308 20402
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13188 19910 13308 19938
rect 13464 19922 13492 20198
rect 13832 19990 13860 20470
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13452 19916 13504 19922
rect 13188 18358 13216 19910
rect 13452 19858 13504 19864
rect 14384 19854 14412 20198
rect 14476 20058 14504 20402
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14752 19922 14780 20402
rect 14844 19990 14872 20402
rect 15396 20398 15424 25230
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15672 23730 15700 25094
rect 15948 23798 15976 25638
rect 16132 25294 16160 25842
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 15764 23050 15792 23666
rect 15752 23044 15804 23050
rect 15752 22986 15804 22992
rect 15764 22778 15792 22986
rect 16132 22982 16160 23666
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 16040 20466 16068 22714
rect 16132 22642 16160 22918
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16132 22094 16160 22578
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 16132 22066 16344 22094
rect 16316 20466 16344 22066
rect 16592 21894 16620 22510
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16684 20602 16712 26522
rect 16776 25974 16804 27542
rect 17144 27334 17172 28018
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 16948 27056 17000 27062
rect 16948 26998 17000 27004
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16764 25968 16816 25974
rect 16764 25910 16816 25916
rect 16868 25906 16896 26930
rect 16960 25974 16988 26998
rect 16948 25968 17000 25974
rect 16948 25910 17000 25916
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16868 24886 16896 25842
rect 17144 25294 17172 27270
rect 17512 27062 17540 28970
rect 17604 28626 17632 33594
rect 17788 33522 17816 34138
rect 18616 34066 18644 34546
rect 18696 34128 18748 34134
rect 18696 34070 18748 34076
rect 18604 34060 18656 34066
rect 18604 34002 18656 34008
rect 18052 33924 18104 33930
rect 18052 33866 18104 33872
rect 17868 33856 17920 33862
rect 17868 33798 17920 33804
rect 18064 33810 18092 33866
rect 17880 33590 17908 33798
rect 18064 33782 18184 33810
rect 18156 33590 18184 33782
rect 17868 33584 17920 33590
rect 17868 33526 17920 33532
rect 18144 33584 18196 33590
rect 18144 33526 18196 33532
rect 17776 33516 17828 33522
rect 17776 33458 17828 33464
rect 17788 29714 17816 33458
rect 18616 32978 18644 34002
rect 18604 32972 18656 32978
rect 18604 32914 18656 32920
rect 18708 32910 18736 34070
rect 18892 33862 18920 34546
rect 19352 34474 19380 34886
rect 19444 34610 19472 35022
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19340 34468 19392 34474
rect 19340 34410 19392 34416
rect 19536 34406 19564 35090
rect 19616 34536 19668 34542
rect 19616 34478 19668 34484
rect 19524 34400 19576 34406
rect 19524 34342 19576 34348
rect 19156 34060 19208 34066
rect 19156 34002 19208 34008
rect 18880 33856 18932 33862
rect 18880 33798 18932 33804
rect 19168 33658 19196 34002
rect 19248 33856 19300 33862
rect 19248 33798 19300 33804
rect 19156 33652 19208 33658
rect 19156 33594 19208 33600
rect 19260 33522 19288 33798
rect 19248 33516 19300 33522
rect 19248 33458 19300 33464
rect 19536 33318 19564 34342
rect 19524 33312 19576 33318
rect 19524 33254 19576 33260
rect 18696 32904 18748 32910
rect 18696 32846 18748 32852
rect 19536 32774 19564 33254
rect 19628 33114 19656 34478
rect 19904 33590 19932 36042
rect 20272 34610 20300 38150
rect 20536 38004 20588 38010
rect 20536 37946 20588 37952
rect 20548 35894 20576 37946
rect 20548 35866 20668 35894
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 20364 34746 20392 35634
rect 20640 34950 20668 35866
rect 20720 35488 20772 35494
rect 20720 35430 20772 35436
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 20352 34740 20404 34746
rect 20352 34682 20404 34688
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 19984 33924 20036 33930
rect 19984 33866 20036 33872
rect 19892 33584 19944 33590
rect 19892 33526 19944 33532
rect 19616 33108 19668 33114
rect 19616 33050 19668 33056
rect 19248 32768 19300 32774
rect 19248 32710 19300 32716
rect 19524 32768 19576 32774
rect 19524 32710 19576 32716
rect 19260 32434 19288 32710
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17776 29708 17828 29714
rect 17776 29650 17828 29656
rect 17592 28620 17644 28626
rect 17592 28562 17644 28568
rect 17604 28506 17632 28562
rect 17880 28558 17908 32166
rect 19340 30184 19392 30190
rect 19340 30126 19392 30132
rect 19352 29170 19380 30126
rect 18328 29164 18380 29170
rect 18328 29106 18380 29112
rect 18420 29164 18472 29170
rect 18420 29106 18472 29112
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 17868 28552 17920 28558
rect 17604 28478 17724 28506
rect 17868 28494 17920 28500
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17604 28082 17632 28358
rect 17696 28150 17724 28478
rect 17684 28144 17736 28150
rect 17684 28086 17736 28092
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 17880 27470 17908 28494
rect 17960 28484 18012 28490
rect 17960 28426 18012 28432
rect 17972 27470 18000 28426
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18156 27606 18184 27950
rect 18248 27674 18276 28494
rect 18340 28218 18368 29106
rect 18432 28762 18460 29106
rect 18420 28756 18472 28762
rect 18420 28698 18472 28704
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 18328 28212 18380 28218
rect 18328 28154 18380 28160
rect 18236 27668 18288 27674
rect 18236 27610 18288 27616
rect 18144 27600 18196 27606
rect 18144 27542 18196 27548
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17500 27056 17552 27062
rect 17500 26998 17552 27004
rect 17604 26042 17632 27406
rect 17684 27396 17736 27402
rect 17684 27338 17736 27344
rect 17696 27130 17724 27338
rect 17684 27124 17736 27130
rect 17684 27066 17736 27072
rect 17972 26994 18000 27406
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 18248 26858 18276 27610
rect 19352 27606 19380 28358
rect 19444 28218 19472 28562
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19432 28212 19484 28218
rect 19432 28154 19484 28160
rect 19616 28076 19668 28082
rect 19616 28018 19668 28024
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 19064 27464 19116 27470
rect 19064 27406 19116 27412
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 17868 26512 17920 26518
rect 17868 26454 17920 26460
rect 17592 26036 17644 26042
rect 17592 25978 17644 25984
rect 17880 25906 17908 26454
rect 18984 26314 19012 27406
rect 19076 27130 19104 27406
rect 19064 27124 19116 27130
rect 19064 27066 19116 27072
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 19260 26382 19288 26930
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19628 26314 19656 28018
rect 19812 27690 19840 28494
rect 19720 27674 19840 27690
rect 19708 27668 19840 27674
rect 19760 27662 19840 27668
rect 19708 27610 19760 27616
rect 19812 26518 19840 27662
rect 19904 26586 19932 33526
rect 19996 32570 20024 33866
rect 20732 33810 20760 35430
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20904 35080 20956 35086
rect 20904 35022 20956 35028
rect 20824 34746 20852 35022
rect 20812 34740 20864 34746
rect 20812 34682 20864 34688
rect 20732 33782 20852 33810
rect 20720 32836 20772 32842
rect 20720 32778 20772 32784
rect 20732 32570 20760 32778
rect 19984 32564 20036 32570
rect 19984 32506 20036 32512
rect 20720 32564 20772 32570
rect 20720 32506 20772 32512
rect 20824 32434 20852 33782
rect 20812 32428 20864 32434
rect 20812 32370 20864 32376
rect 20916 31958 20944 35022
rect 20996 34944 21048 34950
rect 20996 34886 21048 34892
rect 21008 33454 21036 34886
rect 21376 34678 21404 39374
rect 22848 37262 22876 41550
rect 23480 41540 23532 41546
rect 23480 41482 23532 41488
rect 23492 41274 23520 41482
rect 24400 41472 24452 41478
rect 24400 41414 24452 41420
rect 23480 41268 23532 41274
rect 23480 41210 23532 41216
rect 23388 41132 23440 41138
rect 23388 41074 23440 41080
rect 24124 41132 24176 41138
rect 24124 41074 24176 41080
rect 23204 41064 23256 41070
rect 23204 41006 23256 41012
rect 23216 40730 23244 41006
rect 23204 40724 23256 40730
rect 23204 40666 23256 40672
rect 23112 40044 23164 40050
rect 23112 39986 23164 39992
rect 23296 40044 23348 40050
rect 23296 39986 23348 39992
rect 23124 39302 23152 39986
rect 23308 39302 23336 39986
rect 23112 39296 23164 39302
rect 23112 39238 23164 39244
rect 23296 39296 23348 39302
rect 23296 39238 23348 39244
rect 23124 38894 23152 39238
rect 23308 38962 23336 39238
rect 23296 38956 23348 38962
rect 23296 38898 23348 38904
rect 23112 38888 23164 38894
rect 23112 38830 23164 38836
rect 23296 37664 23348 37670
rect 23296 37606 23348 37612
rect 22836 37256 22888 37262
rect 22836 37198 22888 37204
rect 22848 36786 22876 37198
rect 23204 37188 23256 37194
rect 23204 37130 23256 37136
rect 23216 36922 23244 37130
rect 23204 36916 23256 36922
rect 23204 36858 23256 36864
rect 23308 36786 23336 37606
rect 23400 36854 23428 41074
rect 23480 40588 23532 40594
rect 23480 40530 23532 40536
rect 23492 40186 23520 40530
rect 24136 40526 24164 41074
rect 24216 40724 24268 40730
rect 24216 40666 24268 40672
rect 24124 40520 24176 40526
rect 24124 40462 24176 40468
rect 23940 40384 23992 40390
rect 23940 40326 23992 40332
rect 23480 40180 23532 40186
rect 23480 40122 23532 40128
rect 23952 40050 23980 40326
rect 23940 40044 23992 40050
rect 23940 39986 23992 39992
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23676 39642 23704 39918
rect 24032 39840 24084 39846
rect 24032 39782 24084 39788
rect 23572 39636 23624 39642
rect 23572 39578 23624 39584
rect 23664 39636 23716 39642
rect 23664 39578 23716 39584
rect 23584 39370 23612 39578
rect 24044 39438 24072 39782
rect 24228 39438 24256 40666
rect 24412 40526 24440 41414
rect 24400 40520 24452 40526
rect 24400 40462 24452 40468
rect 24308 40384 24360 40390
rect 24308 40326 24360 40332
rect 24032 39432 24084 39438
rect 24032 39374 24084 39380
rect 24216 39432 24268 39438
rect 24216 39374 24268 39380
rect 23572 39364 23624 39370
rect 23572 39306 23624 39312
rect 23572 38820 23624 38826
rect 23572 38762 23624 38768
rect 23584 38010 23612 38762
rect 23572 38004 23624 38010
rect 23572 37946 23624 37952
rect 23664 37868 23716 37874
rect 23664 37810 23716 37816
rect 23676 37482 23704 37810
rect 23676 37466 23796 37482
rect 23676 37460 23808 37466
rect 23676 37454 23756 37460
rect 23388 36848 23440 36854
rect 23388 36790 23440 36796
rect 22836 36780 22888 36786
rect 22836 36722 22888 36728
rect 23296 36780 23348 36786
rect 23296 36722 23348 36728
rect 22848 36242 22876 36722
rect 22836 36236 22888 36242
rect 22836 36178 22888 36184
rect 22008 35012 22060 35018
rect 22008 34954 22060 34960
rect 21364 34672 21416 34678
rect 21364 34614 21416 34620
rect 22020 34610 22048 34954
rect 22928 34672 22980 34678
rect 22928 34614 22980 34620
rect 22008 34604 22060 34610
rect 22008 34546 22060 34552
rect 22100 34536 22152 34542
rect 22100 34478 22152 34484
rect 22112 34066 22140 34478
rect 22940 34474 22968 34614
rect 23676 34610 23704 37454
rect 23756 37402 23808 37408
rect 24044 37126 24072 39374
rect 24032 37120 24084 37126
rect 24032 37062 24084 37068
rect 24320 34678 24348 40326
rect 24412 40050 24440 40462
rect 24400 40044 24452 40050
rect 24400 39986 24452 39992
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 24412 37126 24440 37198
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24308 34672 24360 34678
rect 24308 34614 24360 34620
rect 23664 34604 23716 34610
rect 23664 34546 23716 34552
rect 22928 34468 22980 34474
rect 22928 34410 22980 34416
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 21180 33992 21232 33998
rect 21180 33934 21232 33940
rect 21272 33992 21324 33998
rect 21272 33934 21324 33940
rect 21192 33658 21220 33934
rect 21180 33652 21232 33658
rect 21180 33594 21232 33600
rect 21192 33454 21220 33594
rect 20996 33448 21048 33454
rect 20996 33390 21048 33396
rect 21180 33448 21232 33454
rect 21180 33390 21232 33396
rect 21008 32434 21036 33390
rect 21192 33046 21220 33390
rect 21284 33318 21312 33934
rect 22940 33930 22968 34410
rect 23204 34196 23256 34202
rect 23204 34138 23256 34144
rect 22468 33924 22520 33930
rect 22468 33866 22520 33872
rect 22928 33924 22980 33930
rect 22928 33866 22980 33872
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22100 33516 22152 33522
rect 22100 33458 22152 33464
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21284 33114 21312 33254
rect 22112 33114 22140 33458
rect 21272 33108 21324 33114
rect 21272 33050 21324 33056
rect 22100 33108 22152 33114
rect 22100 33050 22152 33056
rect 21180 33040 21232 33046
rect 21180 32982 21232 32988
rect 20996 32428 21048 32434
rect 20996 32370 21048 32376
rect 20904 31952 20956 31958
rect 20904 31894 20956 31900
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19996 28558 20024 29106
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 20904 28552 20956 28558
rect 20904 28494 20956 28500
rect 20260 28484 20312 28490
rect 20260 28426 20312 28432
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 19996 26994 20024 27270
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19996 26586 20024 26930
rect 19892 26580 19944 26586
rect 19892 26522 19944 26528
rect 19984 26580 20036 26586
rect 19984 26522 20036 26528
rect 19800 26512 19852 26518
rect 19800 26454 19852 26460
rect 20272 26382 20300 28426
rect 20812 28416 20864 28422
rect 20812 28358 20864 28364
rect 20824 27470 20852 28358
rect 20916 27674 20944 28494
rect 21192 28082 21220 32982
rect 21284 32502 21312 33050
rect 21824 32972 21876 32978
rect 21824 32914 21876 32920
rect 21836 32502 21864 32914
rect 22192 32836 22244 32842
rect 22192 32778 22244 32784
rect 22204 32570 22232 32778
rect 22296 32774 22324 33798
rect 22480 33522 22508 33866
rect 22468 33516 22520 33522
rect 22468 33458 22520 33464
rect 22376 32836 22428 32842
rect 22376 32778 22428 32784
rect 22284 32768 22336 32774
rect 22284 32710 22336 32716
rect 22192 32564 22244 32570
rect 22192 32506 22244 32512
rect 21272 32496 21324 32502
rect 21272 32438 21324 32444
rect 21824 32496 21876 32502
rect 21824 32438 21876 32444
rect 22388 32434 22416 32778
rect 22480 32434 22508 33458
rect 22940 33114 22968 33866
rect 23216 33658 23244 34138
rect 24032 33856 24084 33862
rect 24032 33798 24084 33804
rect 23204 33652 23256 33658
rect 23204 33594 23256 33600
rect 23296 33312 23348 33318
rect 23296 33254 23348 33260
rect 22928 33108 22980 33114
rect 22928 33050 22980 33056
rect 23308 32910 23336 33254
rect 24044 32910 24072 33798
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 24032 32904 24084 32910
rect 24032 32846 24084 32852
rect 24308 32904 24360 32910
rect 24308 32846 24360 32852
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 24216 32768 24268 32774
rect 24216 32710 24268 32716
rect 23308 32434 23336 32710
rect 22376 32428 22428 32434
rect 22376 32370 22428 32376
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 21272 31952 21324 31958
rect 21272 31894 21324 31900
rect 21284 28558 21312 31894
rect 24228 31822 24256 32710
rect 24320 31958 24348 32846
rect 24400 32428 24452 32434
rect 24400 32370 24452 32376
rect 24412 32026 24440 32370
rect 24400 32020 24452 32026
rect 24400 31962 24452 31968
rect 24308 31952 24360 31958
rect 24308 31894 24360 31900
rect 24216 31816 24268 31822
rect 24216 31758 24268 31764
rect 22376 28688 22428 28694
rect 22376 28630 22428 28636
rect 21272 28552 21324 28558
rect 21272 28494 21324 28500
rect 22008 28144 22060 28150
rect 22008 28086 22060 28092
rect 21180 28076 21232 28082
rect 21180 28018 21232 28024
rect 20904 27668 20956 27674
rect 20904 27610 20956 27616
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20824 26790 20852 27406
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20916 26382 20944 27610
rect 21192 27402 21220 28018
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 21560 27538 21588 27814
rect 22020 27538 22048 28086
rect 21548 27532 21600 27538
rect 21548 27474 21600 27480
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 22388 27470 22416 28630
rect 21824 27464 21876 27470
rect 21824 27406 21876 27412
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 21548 27396 21600 27402
rect 21548 27338 21600 27344
rect 21192 26994 21220 27338
rect 21560 27062 21588 27338
rect 21548 27056 21600 27062
rect 21548 26998 21600 27004
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 21836 26586 21864 27406
rect 21824 26580 21876 26586
rect 21824 26522 21876 26528
rect 24504 26450 24532 45526
rect 26516 41608 26568 41614
rect 26516 41550 26568 41556
rect 26792 41608 26844 41614
rect 26792 41550 26844 41556
rect 26424 41132 26476 41138
rect 26424 41074 26476 41080
rect 24584 41064 24636 41070
rect 24584 41006 24636 41012
rect 26148 41064 26200 41070
rect 26148 41006 26200 41012
rect 24596 37738 24624 41006
rect 26160 40474 26188 41006
rect 26332 40520 26384 40526
rect 26330 40488 26332 40497
rect 26384 40488 26386 40497
rect 26160 40458 26280 40474
rect 26160 40452 26292 40458
rect 26160 40446 26240 40452
rect 26160 40186 26188 40446
rect 26330 40423 26386 40432
rect 26240 40394 26292 40400
rect 26436 40186 26464 41074
rect 26148 40180 26200 40186
rect 26148 40122 26200 40128
rect 26424 40180 26476 40186
rect 26424 40122 26476 40128
rect 24676 40044 24728 40050
rect 24676 39986 24728 39992
rect 26240 40044 26292 40050
rect 26240 39986 26292 39992
rect 24688 39574 24716 39986
rect 24676 39568 24728 39574
rect 24676 39510 24728 39516
rect 26252 37806 26280 39986
rect 26240 37800 26292 37806
rect 26240 37742 26292 37748
rect 24584 37732 24636 37738
rect 24584 37674 24636 37680
rect 26528 37262 26556 41550
rect 26700 41472 26752 41478
rect 26700 41414 26752 41420
rect 26712 41206 26740 41414
rect 26700 41200 26752 41206
rect 26700 41142 26752 41148
rect 26804 40730 26832 41550
rect 26976 41064 27028 41070
rect 26976 41006 27028 41012
rect 26608 40724 26660 40730
rect 26792 40724 26844 40730
rect 26660 40684 26740 40712
rect 26608 40666 26660 40672
rect 26712 40594 26740 40684
rect 26792 40666 26844 40672
rect 26700 40588 26752 40594
rect 26700 40530 26752 40536
rect 26712 40050 26740 40530
rect 26700 40044 26752 40050
rect 26700 39986 26752 39992
rect 26884 38548 26936 38554
rect 26884 38490 26936 38496
rect 26896 37738 26924 38490
rect 26884 37732 26936 37738
rect 26884 37674 26936 37680
rect 26896 37262 26924 37674
rect 26516 37256 26568 37262
rect 26516 37198 26568 37204
rect 26884 37256 26936 37262
rect 26884 37198 26936 37204
rect 26528 35170 26556 37198
rect 26608 37188 26660 37194
rect 26608 37130 26660 37136
rect 26620 36854 26648 37130
rect 26884 37120 26936 37126
rect 26988 37074 27016 41006
rect 27160 40928 27212 40934
rect 27160 40870 27212 40876
rect 27712 40928 27764 40934
rect 27712 40870 27764 40876
rect 27172 40594 27200 40870
rect 27160 40588 27212 40594
rect 27160 40530 27212 40536
rect 27344 40588 27396 40594
rect 27344 40530 27396 40536
rect 27252 40384 27304 40390
rect 27252 40326 27304 40332
rect 27160 38412 27212 38418
rect 27160 38354 27212 38360
rect 27068 38208 27120 38214
rect 27068 38150 27120 38156
rect 27080 37262 27108 38150
rect 27172 38010 27200 38354
rect 27160 38004 27212 38010
rect 27160 37946 27212 37952
rect 27160 37868 27212 37874
rect 27160 37810 27212 37816
rect 27172 37262 27200 37810
rect 27068 37256 27120 37262
rect 27068 37198 27120 37204
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 26936 37068 27016 37074
rect 26884 37062 27016 37068
rect 26896 37046 27016 37062
rect 26608 36848 26660 36854
rect 26608 36790 26660 36796
rect 26988 36786 27016 37046
rect 26976 36780 27028 36786
rect 26976 36722 27028 36728
rect 26792 35624 26844 35630
rect 26792 35566 26844 35572
rect 26528 35142 26648 35170
rect 25228 34740 25280 34746
rect 25228 34682 25280 34688
rect 24860 34536 24912 34542
rect 24860 34478 24912 34484
rect 24872 33114 24900 34478
rect 25240 33998 25268 34682
rect 26516 34604 26568 34610
rect 26516 34546 26568 34552
rect 25596 34536 25648 34542
rect 25596 34478 25648 34484
rect 25412 34400 25464 34406
rect 25412 34342 25464 34348
rect 25424 33998 25452 34342
rect 25608 33998 25636 34478
rect 25228 33992 25280 33998
rect 25228 33934 25280 33940
rect 25412 33992 25464 33998
rect 25412 33934 25464 33940
rect 25596 33992 25648 33998
rect 25596 33934 25648 33940
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24872 32978 24900 33050
rect 24860 32972 24912 32978
rect 24860 32914 24912 32920
rect 24768 32768 24820 32774
rect 24768 32710 24820 32716
rect 24780 32026 24808 32710
rect 24872 32570 24900 32914
rect 25608 32842 25636 33934
rect 26528 33862 26556 34546
rect 26620 34474 26648 35142
rect 26804 34678 26832 35566
rect 26988 35086 27016 36722
rect 26976 35080 27028 35086
rect 26976 35022 27028 35028
rect 26792 34672 26844 34678
rect 26792 34614 26844 34620
rect 26976 34604 27028 34610
rect 26976 34546 27028 34552
rect 26608 34468 26660 34474
rect 26608 34410 26660 34416
rect 26516 33856 26568 33862
rect 26516 33798 26568 33804
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 25596 32836 25648 32842
rect 25596 32778 25648 32784
rect 25688 32836 25740 32842
rect 25688 32778 25740 32784
rect 25608 32570 25636 32778
rect 24860 32564 24912 32570
rect 24860 32506 24912 32512
rect 25596 32564 25648 32570
rect 25596 32506 25648 32512
rect 24768 32020 24820 32026
rect 24768 31962 24820 31968
rect 24872 31958 24900 32506
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 24860 31952 24912 31958
rect 24860 31894 24912 31900
rect 25044 31748 25096 31754
rect 25044 31690 25096 31696
rect 24952 31680 25004 31686
rect 24952 31622 25004 31628
rect 24964 31346 24992 31622
rect 25056 31346 25084 31690
rect 25424 31482 25452 32370
rect 25700 31822 25728 32778
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 26068 31890 26096 32506
rect 26160 32026 26188 32846
rect 26148 32020 26200 32026
rect 26148 31962 26200 31968
rect 26056 31884 26108 31890
rect 26056 31826 26108 31832
rect 25688 31816 25740 31822
rect 25688 31758 25740 31764
rect 25412 31476 25464 31482
rect 25412 31418 25464 31424
rect 25700 31346 25728 31758
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 25688 31340 25740 31346
rect 25688 31282 25740 31288
rect 26160 31278 26188 31962
rect 26528 31890 26556 33798
rect 26620 33522 26648 34410
rect 26988 34202 27016 34546
rect 27264 34542 27292 40326
rect 27356 38554 27384 40530
rect 27436 40520 27488 40526
rect 27724 40497 27752 40870
rect 27436 40462 27488 40468
rect 27710 40488 27766 40497
rect 27448 40118 27476 40462
rect 27710 40423 27766 40432
rect 27528 40384 27580 40390
rect 27528 40326 27580 40332
rect 27436 40112 27488 40118
rect 27436 40054 27488 40060
rect 27344 38548 27396 38554
rect 27344 38490 27396 38496
rect 27540 38350 27568 40326
rect 27724 40118 27752 40423
rect 27896 40384 27948 40390
rect 27896 40326 27948 40332
rect 27908 40186 27936 40326
rect 27896 40180 27948 40186
rect 27896 40122 27948 40128
rect 27712 40112 27764 40118
rect 27712 40054 27764 40060
rect 27908 39914 27936 40122
rect 27896 39908 27948 39914
rect 27896 39850 27948 39856
rect 27528 38344 27580 38350
rect 27528 38286 27580 38292
rect 27344 37868 27396 37874
rect 27344 37810 27396 37816
rect 27356 36922 27384 37810
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 27344 36916 27396 36922
rect 27344 36858 27396 36864
rect 27356 34746 27384 36858
rect 28460 36582 28488 37198
rect 28448 36576 28500 36582
rect 28448 36518 28500 36524
rect 28264 35692 28316 35698
rect 28264 35634 28316 35640
rect 27620 35488 27672 35494
rect 27620 35430 27672 35436
rect 27632 35086 27660 35430
rect 28276 35290 28304 35634
rect 28448 35488 28500 35494
rect 28446 35456 28448 35465
rect 28500 35456 28502 35465
rect 28446 35391 28502 35400
rect 28264 35284 28316 35290
rect 28264 35226 28316 35232
rect 27620 35080 27672 35086
rect 27620 35022 27672 35028
rect 27344 34740 27396 34746
rect 27344 34682 27396 34688
rect 27356 34592 27384 34682
rect 27436 34604 27488 34610
rect 27356 34564 27436 34592
rect 27436 34546 27488 34552
rect 27252 34536 27304 34542
rect 27252 34478 27304 34484
rect 27988 34536 28040 34542
rect 27988 34478 28040 34484
rect 26976 34196 27028 34202
rect 26976 34138 27028 34144
rect 27264 33930 27292 34478
rect 28000 34066 28028 34478
rect 27988 34060 28040 34066
rect 27988 34002 28040 34008
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 26608 33516 26660 33522
rect 26608 33458 26660 33464
rect 26620 32994 26648 33458
rect 26620 32966 26832 32994
rect 28000 32978 28028 34002
rect 26804 32910 26832 32966
rect 27988 32972 28040 32978
rect 27988 32914 28040 32920
rect 26792 32904 26844 32910
rect 26844 32852 26924 32858
rect 26792 32846 26924 32852
rect 26804 32830 26924 32846
rect 26792 32768 26844 32774
rect 26792 32710 26844 32716
rect 26516 31884 26568 31890
rect 26516 31826 26568 31832
rect 26804 31822 26832 32710
rect 26792 31816 26844 31822
rect 26792 31758 26844 31764
rect 26148 31272 26200 31278
rect 26148 31214 26200 31220
rect 24492 26444 24544 26450
rect 24492 26386 24544 26392
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 18972 26308 19024 26314
rect 18972 26250 19024 26256
rect 19616 26308 19668 26314
rect 19616 26250 19668 26256
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 16856 24880 16908 24886
rect 16856 24822 16908 24828
rect 17236 23866 17264 25842
rect 18984 23866 19012 26250
rect 26896 26234 26924 32830
rect 28000 32570 28028 32914
rect 27988 32564 28040 32570
rect 27988 32506 28040 32512
rect 26976 32428 27028 32434
rect 26976 32370 27028 32376
rect 27068 32428 27120 32434
rect 27068 32370 27120 32376
rect 26988 30258 27016 32370
rect 27080 32026 27108 32370
rect 27068 32020 27120 32026
rect 27068 31962 27120 31968
rect 28448 31952 28500 31958
rect 28448 31894 28500 31900
rect 28356 31816 28408 31822
rect 28356 31758 28408 31764
rect 26976 30252 27028 30258
rect 26976 30194 27028 30200
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 27080 29034 27108 30194
rect 28368 30122 28396 31758
rect 28460 31385 28488 31894
rect 28446 31376 28502 31385
rect 28446 31311 28502 31320
rect 28356 30116 28408 30122
rect 28356 30058 28408 30064
rect 27068 29028 27120 29034
rect 27068 28970 27120 28976
rect 28538 27976 28594 27985
rect 28538 27911 28540 27920
rect 28592 27911 28594 27920
rect 28540 27882 28592 27888
rect 26804 26206 26924 26234
rect 19432 25764 19484 25770
rect 19432 25706 19484 25712
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 18972 23860 19024 23866
rect 18972 23802 19024 23808
rect 18144 23792 18196 23798
rect 18144 23734 18196 23740
rect 17960 23656 18012 23662
rect 17960 23598 18012 23604
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16868 23322 16896 23462
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16776 22506 16804 22986
rect 16868 22642 16896 23258
rect 17972 23186 18000 23598
rect 18156 23254 18184 23734
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 18144 23248 18196 23254
rect 18144 23190 18196 23196
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 17144 22030 17172 22918
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 14832 19984 14884 19990
rect 14832 19926 14884 19932
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12912 10810 12940 11018
rect 13188 10810 13216 18294
rect 14752 17678 14780 19858
rect 15396 19854 15424 20334
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15660 19780 15712 19786
rect 15660 19722 15712 19728
rect 15672 19514 15700 19722
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15856 19378 15884 20198
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15948 18222 15976 20402
rect 16040 19530 16068 20402
rect 16316 20058 16344 20402
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 16040 19502 16160 19530
rect 16132 19378 16160 19502
rect 16684 19378 16712 20538
rect 17420 20534 17448 21966
rect 17972 21962 18000 22578
rect 18064 22030 18092 22578
rect 18156 22574 18184 23190
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 18512 22976 18564 22982
rect 18512 22918 18564 22924
rect 18524 22642 18552 22918
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18156 22234 18184 22510
rect 18892 22234 18920 23054
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18880 22228 18932 22234
rect 18880 22170 18932 22176
rect 18616 22030 18644 22170
rect 18892 22094 18920 22170
rect 18800 22066 18920 22094
rect 18800 22030 18828 22066
rect 18984 22030 19012 23598
rect 19444 23526 19472 25706
rect 19616 24880 19668 24886
rect 19616 24822 19668 24828
rect 19628 23798 19656 24822
rect 19616 23792 19668 23798
rect 19616 23734 19668 23740
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19444 23118 19472 23462
rect 19628 23254 19656 23734
rect 19708 23520 19760 23526
rect 19708 23462 19760 23468
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19260 22778 19288 22918
rect 19444 22778 19472 23054
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19444 22098 19472 22714
rect 19628 22506 19656 23190
rect 19720 23050 19748 23462
rect 19708 23044 19760 23050
rect 19708 22986 19760 22992
rect 19616 22500 19668 22506
rect 19616 22442 19668 22448
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 17960 21956 18012 21962
rect 17960 21898 18012 21904
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 17408 20528 17460 20534
rect 17408 20470 17460 20476
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16776 19446 16804 19654
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 16132 18290 16160 19314
rect 17972 18290 18000 19314
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 15212 17610 15240 18022
rect 16132 17882 16160 18226
rect 18524 18222 18552 21830
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 19260 18290 19288 18702
rect 19616 18692 19668 18698
rect 19616 18634 19668 18640
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 18340 17678 18368 18022
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 18340 17202 18368 17614
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16868 16590 16896 16934
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17328 15910 17356 16526
rect 18156 16182 18184 17070
rect 18248 16454 18276 17070
rect 18340 16794 18368 17138
rect 18432 16794 18460 17614
rect 18524 17610 18552 18158
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 18248 16250 18276 16390
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 13740 15094 13768 15846
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13372 14346 13400 14486
rect 13464 14414 13492 14962
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13372 13530 13400 14282
rect 13452 14272 13504 14278
rect 13556 14226 13584 14894
rect 13648 14550 13676 14962
rect 13740 14618 13768 15030
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13740 14362 13768 14554
rect 14936 14550 14964 14962
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 13648 14346 13768 14362
rect 13636 14340 13768 14346
rect 13688 14334 13768 14340
rect 15476 14340 15528 14346
rect 13636 14282 13688 14288
rect 15476 14282 15528 14288
rect 13504 14220 13584 14226
rect 13452 14214 13584 14220
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 13464 14198 13584 14214
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13464 12238 13492 14198
rect 15304 13326 15332 14214
rect 15488 13530 15516 14282
rect 16224 13938 16252 14758
rect 17236 14414 17264 15030
rect 17328 15026 17356 15846
rect 17788 15706 17816 16050
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18156 15706 18184 15846
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18248 15502 18276 16186
rect 18340 16114 18368 16730
rect 18512 16516 18564 16522
rect 18512 16458 18564 16464
rect 18524 16250 18552 16458
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17328 14414 17356 14962
rect 18248 14482 18276 15438
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18340 14414 18368 14758
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15488 13326 15516 13466
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 13190 15516 13262
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16040 12918 16068 13126
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16132 12850 16160 13126
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 13464 11354 13492 12174
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 15120 11218 15148 11494
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15212 11150 15240 12174
rect 16132 11830 16160 12786
rect 16224 11830 16252 13874
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16592 11898 16620 13194
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15488 11354 15516 11698
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15212 10826 15240 11086
rect 15764 11082 15792 11698
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16040 11218 16068 11562
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 13176 10804 13228 10810
rect 15212 10798 15332 10826
rect 13176 10746 13228 10752
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11532 9722 11560 9862
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10520 9042 10640 9058
rect 10520 9036 10652 9042
rect 10520 9030 10600 9036
rect 10600 8978 10652 8984
rect 10796 8974 10824 9386
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10428 8634 10456 8842
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10980 8498 11008 8978
rect 11164 8498 11192 9318
rect 12176 9178 12204 9522
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 12360 8430 12388 8842
rect 13188 8566 13216 10746
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14476 10062 14504 10542
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14476 9518 14504 9998
rect 14568 9654 14596 10678
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15212 10266 15240 10610
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 15028 9654 15056 9998
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15200 9648 15252 9654
rect 15304 9636 15332 10798
rect 15488 10062 15516 10950
rect 15764 10810 15792 11018
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 16040 9722 16068 11154
rect 16500 11150 16528 11630
rect 16592 11286 16620 11834
rect 16776 11830 16804 13330
rect 16960 12782 16988 14350
rect 17236 13818 17264 14350
rect 17052 13790 17264 13818
rect 17052 13258 17080 13790
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17236 13326 17264 13670
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16960 12442 16988 12718
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 17972 10674 18000 12650
rect 18432 11762 18460 14350
rect 18708 14006 18736 18226
rect 19260 18086 19288 18226
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19628 17882 19656 18634
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18800 17270 18828 17478
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18892 16726 18920 17614
rect 20180 17542 20208 17614
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20456 17338 20484 18226
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20732 17202 20760 18634
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20824 17270 20852 17682
rect 20916 17678 20944 18702
rect 21100 18630 21128 18770
rect 22112 18766 22140 18838
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 21100 17678 21128 18566
rect 21192 17814 21220 18702
rect 21468 17814 21496 18702
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21180 17808 21232 17814
rect 21180 17750 21232 17756
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19720 16794 19748 17002
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19168 15570 19196 15846
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19352 14618 19380 15370
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19444 14498 19472 15302
rect 19720 14550 19748 16730
rect 19812 16590 19840 16934
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 20640 15502 20668 16934
rect 20824 15502 20852 17206
rect 20916 17202 20944 17614
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 21008 17202 21036 17478
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21100 16998 21128 17614
rect 21192 17338 21220 17750
rect 21468 17338 21496 17750
rect 21560 17746 21588 18022
rect 21548 17740 21600 17746
rect 21548 17682 21600 17688
rect 22112 17610 22140 18702
rect 23664 18692 23716 18698
rect 23664 18634 23716 18640
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22296 17882 22324 18226
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 22112 17202 22140 17546
rect 22572 17338 22600 17614
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 23124 17202 23152 18566
rect 23492 17202 23520 18566
rect 23676 18426 23704 18634
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23676 17746 23704 18362
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 23676 16574 23704 17682
rect 23768 17338 23796 18226
rect 23952 17882 23980 18702
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24044 17746 24072 17818
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 24308 17604 24360 17610
rect 24308 17546 24360 17552
rect 23756 17332 23808 17338
rect 23756 17274 23808 17280
rect 23492 16546 23704 16574
rect 21456 16176 21508 16182
rect 21456 16118 21508 16124
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 19904 14550 19932 15438
rect 19996 14618 20024 15438
rect 20260 15428 20312 15434
rect 20260 15370 20312 15376
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19352 14482 19472 14498
rect 19708 14544 19760 14550
rect 19708 14486 19760 14492
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19340 14476 19472 14482
rect 19392 14470 19472 14476
rect 19340 14418 19392 14424
rect 19720 14414 19748 14486
rect 20272 14482 20300 15370
rect 20824 14550 20852 15438
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18052 11620 18104 11626
rect 18052 11562 18104 11568
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 18064 10606 18092 11562
rect 18432 10962 18460 11698
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18340 10934 18460 10962
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 15252 9608 15332 9636
rect 15200 9590 15252 9596
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14280 8968 14332 8974
rect 14476 8956 14504 9454
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14332 8928 14504 8956
rect 14280 8910 14332 8916
rect 14476 8566 14504 8928
rect 14740 8900 14792 8906
rect 14740 8842 14792 8848
rect 14752 8634 14780 8842
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14936 8498 14964 9318
rect 15028 8974 15056 9590
rect 15304 9178 15332 9608
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 15304 8498 15332 9114
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15396 8430 15424 9522
rect 17972 8974 18000 9862
rect 18064 9586 18092 10542
rect 18156 10062 18184 10542
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9722 18184 9862
rect 18248 9722 18276 10610
rect 18340 10062 18368 10934
rect 18800 10606 18828 11630
rect 18892 10674 18920 14350
rect 21468 13326 21496 16118
rect 23492 16114 23520 16546
rect 24320 16114 24348 17546
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24412 17270 24440 17478
rect 24780 17270 24808 17750
rect 24872 17610 24900 18022
rect 25240 17882 25268 18226
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25412 17672 25464 17678
rect 25412 17614 25464 17620
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24400 17264 24452 17270
rect 24400 17206 24452 17212
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 25424 17066 25452 17614
rect 25516 17202 25544 18634
rect 26240 18080 26292 18086
rect 26240 18022 26292 18028
rect 26516 18080 26568 18086
rect 26516 18022 26568 18028
rect 25872 17740 25924 17746
rect 25872 17682 25924 17688
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25608 17338 25636 17478
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25516 17082 25544 17138
rect 25412 17060 25464 17066
rect 25516 17054 25636 17082
rect 25412 17002 25464 17008
rect 25608 16794 25636 17054
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 25608 16674 25636 16730
rect 25424 16646 25636 16674
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24872 16114 24900 16390
rect 23296 16108 23348 16114
rect 23296 16050 23348 16056
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21560 14346 21588 15438
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 21744 15026 21772 15302
rect 22112 15094 22140 15302
rect 22204 15094 22232 15982
rect 23308 15162 23336 16050
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 19536 10606 19564 10746
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 18800 10470 18828 10542
rect 19340 10532 19392 10538
rect 19340 10474 19392 10480
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 18432 10130 18460 10406
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18524 9926 18552 10066
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18616 9586 18644 9930
rect 19076 9586 19104 9998
rect 19168 9586 19196 10406
rect 19352 10130 19380 10474
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19352 9654 19380 9930
rect 19444 9722 19472 10542
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8498 17264 8774
rect 18708 8498 18736 8842
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18892 8498 18920 8774
rect 19076 8634 19104 9522
rect 19536 9110 19564 9862
rect 19524 9104 19576 9110
rect 19524 9046 19576 9052
rect 19628 8974 19656 10678
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19720 9042 19748 9862
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 20088 8974 20116 9454
rect 20732 9450 20760 13262
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 21192 9518 21220 11766
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21284 10810 21312 11154
rect 21376 11150 21404 12718
rect 21560 12374 21588 14282
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21640 12708 21692 12714
rect 21640 12650 21692 12656
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21468 11354 21496 12242
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21376 10470 21404 11086
rect 21560 11082 21588 12310
rect 21652 12238 21680 12650
rect 21744 12442 21772 13262
rect 21836 12850 21864 13330
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 22020 12918 22048 13126
rect 23400 12986 23428 15982
rect 23492 15026 23520 16050
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 24860 13728 24912 13734
rect 24860 13670 24912 13676
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 24872 13326 24900 13670
rect 25056 13530 25084 13670
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21652 11286 21680 12174
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21376 10198 21404 10406
rect 21364 10192 21416 10198
rect 21364 10134 21416 10140
rect 21560 9586 21588 11018
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 20076 8968 20128 8974
rect 20128 8928 20208 8956
rect 20076 8910 20128 8916
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 10796 7818 10824 8230
rect 19260 7954 19288 8434
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19352 7886 19380 8298
rect 20180 8090 20208 8928
rect 20732 8430 20760 9386
rect 21560 9042 21588 9522
rect 21836 9042 21864 12786
rect 22388 12442 22416 12786
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21928 9518 21956 11154
rect 22296 11150 22324 12174
rect 22388 12102 22416 12378
rect 23308 12306 23336 12786
rect 23400 12442 23428 12922
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 24504 12238 24532 13262
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 24492 12232 24544 12238
rect 24544 12192 24624 12220
rect 24492 12174 24544 12180
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 23032 11830 23060 12174
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 24492 11212 24544 11218
rect 24492 11154 24544 11160
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22008 11076 22060 11082
rect 22008 11018 22060 11024
rect 22020 9586 22048 11018
rect 24504 10674 24532 11154
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24504 10130 24532 10610
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24596 9586 24624 12192
rect 24872 10674 24900 12718
rect 25136 10736 25188 10742
rect 25136 10678 25188 10684
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24780 10266 24808 10610
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24872 10198 24900 10610
rect 25148 10198 25176 10678
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 25136 10192 25188 10198
rect 25136 10134 25188 10140
rect 25240 9926 25268 15846
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25332 12986 25360 13874
rect 25424 13870 25452 16646
rect 25884 16590 25912 17682
rect 26252 16658 26280 18022
rect 26528 17678 26556 18022
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25872 16584 25924 16590
rect 25872 16526 25924 16532
rect 25516 16250 25544 16526
rect 25596 16448 25648 16454
rect 25596 16390 25648 16396
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25608 14074 25636 16390
rect 26528 15978 26556 17614
rect 26516 15972 26568 15978
rect 26516 15914 26568 15920
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 25228 9920 25280 9926
rect 25228 9862 25280 9868
rect 24964 9722 24992 9862
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 25240 9586 25268 9862
rect 25424 9654 25452 13806
rect 25608 12986 25636 14010
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 25700 13530 25728 13874
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25608 10810 25636 12786
rect 25596 10804 25648 10810
rect 25596 10746 25648 10752
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 25608 9654 25636 10202
rect 25976 10062 26004 10610
rect 26804 10266 26832 26206
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 28276 23322 28304 23666
rect 28448 23520 28500 23526
rect 28448 23462 28500 23468
rect 28264 23316 28316 23322
rect 28264 23258 28316 23264
rect 28460 23225 28488 23462
rect 28446 23216 28502 23225
rect 28446 23151 28502 23160
rect 27528 23112 27580 23118
rect 27528 23054 27580 23060
rect 27540 18698 27568 23054
rect 28540 22568 28592 22574
rect 28538 22536 28540 22545
rect 28592 22536 28594 22545
rect 28538 22471 28594 22480
rect 28540 19848 28592 19854
rect 28538 19816 28540 19825
rect 28592 19816 28594 19825
rect 28538 19751 28594 19760
rect 27528 18692 27580 18698
rect 27528 18634 27580 18640
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 28446 16416 28502 16425
rect 28276 16114 28304 16390
rect 28446 16351 28502 16360
rect 28460 16250 28488 16351
rect 28448 16244 28500 16250
rect 28448 16186 28500 16192
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28184 15745 28212 15846
rect 28170 15736 28226 15745
rect 28170 15671 28226 15680
rect 26792 10260 26844 10266
rect 26792 10202 26844 10208
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25596 9648 25648 9654
rect 25596 9590 25648 9596
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21548 9036 21600 9042
rect 21548 8978 21600 8984
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21560 8634 21588 8978
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21836 8498 21864 8978
rect 21928 8974 21956 9046
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 22020 8906 22048 9386
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22008 8900 22060 8906
rect 22008 8842 22060 8848
rect 22388 8838 22416 9114
rect 22480 8974 22508 9318
rect 23952 8974 23980 9318
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 24596 8838 24624 9522
rect 25976 9178 26004 9998
rect 28356 9988 28408 9994
rect 28356 9930 28408 9936
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 22112 8566 22140 8774
rect 28368 8634 28396 9930
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 28540 8492 28592 8498
rect 28540 8434 28592 8440
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 28552 8265 28580 8434
rect 28538 8256 28594 8265
rect 28538 8191 28594 8200
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1306 5304 2382
rect 5184 1278 5304 1306
rect 5184 800 5212 1278
rect 27080 800 27108 2382
rect 5170 0 5226 800
rect 27066 0 27122 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 846 32852 848 32872
rect 848 32852 900 32872
rect 900 32852 902 32872
rect 846 32816 902 32852
rect 846 32172 848 32192
rect 848 32172 900 32192
rect 900 32172 902 32192
rect 846 32136 902 32172
rect 846 31456 902 31512
rect 846 30796 902 30832
rect 846 30776 848 30796
rect 848 30776 900 30796
rect 900 30776 902 30796
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 846 29416 902 29472
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 846 28736 902 28792
rect 12714 31592 12770 31648
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 846 24656 902 24712
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 846 15816 902 15872
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 938 9560 994 9616
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 13542 31592 13598 31648
rect 26330 40468 26332 40488
rect 26332 40468 26384 40488
rect 26384 40468 26386 40488
rect 26330 40432 26386 40468
rect 27710 40432 27766 40488
rect 28446 35436 28448 35456
rect 28448 35436 28500 35456
rect 28500 35436 28502 35456
rect 28446 35400 28502 35436
rect 28446 31320 28502 31376
rect 28538 27940 28594 27976
rect 28538 27920 28540 27940
rect 28540 27920 28592 27940
rect 28592 27920 28594 27940
rect 28446 23160 28502 23216
rect 28538 22516 28540 22536
rect 28540 22516 28592 22536
rect 28592 22516 28594 22536
rect 28538 22480 28594 22516
rect 28538 19796 28540 19816
rect 28540 19796 28592 19816
rect 28592 19796 28594 19816
rect 28538 19760 28594 19796
rect 28446 16360 28502 16416
rect 28170 15680 28226 15736
rect 28538 8200 28594 8256
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 26325 40490 26391 40493
rect 27705 40490 27771 40493
rect 26325 40488 27771 40490
rect 26325 40432 26330 40488
rect 26386 40432 27710 40488
rect 27766 40432 27771 40488
rect 26325 40430 27771 40432
rect 26325 40427 26391 40430
rect 27705 40427 27771 40430
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 28441 35458 28507 35461
rect 29200 35458 30000 35488
rect 28441 35456 30000 35458
rect 28441 35400 28446 35456
rect 28502 35400 30000 35456
rect 28441 35398 30000 35400
rect 28441 35395 28507 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 29200 35368 30000 35398
rect 4210 35327 4526 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 841 32874 907 32877
rect 798 32872 907 32874
rect 798 32816 846 32872
rect 902 32816 907 32872
rect 798 32811 907 32816
rect 798 32768 858 32811
rect 0 32678 858 32768
rect 0 32648 800 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 841 32194 907 32197
rect 798 32192 907 32194
rect 798 32136 846 32192
rect 902 32136 907 32192
rect 798 32131 907 32136
rect 798 32088 858 32131
rect 0 31998 858 32088
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 0 31968 800 31998
rect 12709 31650 12775 31653
rect 13537 31650 13603 31653
rect 12709 31648 13603 31650
rect 12709 31592 12714 31648
rect 12770 31592 13542 31648
rect 13598 31592 13603 31648
rect 12709 31590 13603 31592
rect 12709 31587 12775 31590
rect 13537 31587 13603 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 841 31514 907 31517
rect 798 31512 907 31514
rect 798 31456 846 31512
rect 902 31456 907 31512
rect 798 31451 907 31456
rect 798 31408 858 31451
rect 0 31318 858 31408
rect 28441 31378 28507 31381
rect 29200 31378 30000 31408
rect 28441 31376 30000 31378
rect 28441 31320 28446 31376
rect 28502 31320 30000 31376
rect 28441 31318 30000 31320
rect 0 31288 800 31318
rect 28441 31315 28507 31318
rect 29200 31288 30000 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 841 30834 907 30837
rect 798 30832 907 30834
rect 798 30776 846 30832
rect 902 30776 907 30832
rect 798 30771 907 30776
rect 798 30728 858 30771
rect 0 30638 858 30728
rect 0 30608 800 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 841 29474 907 29477
rect 798 29472 907 29474
rect 798 29416 846 29472
rect 902 29416 907 29472
rect 798 29411 907 29416
rect 798 29368 858 29411
rect 0 29278 858 29368
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 0 29248 800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 841 28794 907 28797
rect 798 28792 907 28794
rect 798 28736 846 28792
rect 902 28736 907 28792
rect 798 28731 907 28736
rect 798 28688 858 28731
rect 0 28598 858 28688
rect 0 28568 800 28598
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 28533 27978 28599 27981
rect 29200 27978 30000 28008
rect 28533 27976 30000 27978
rect 28533 27920 28538 27976
rect 28594 27920 30000 27976
rect 28533 27918 30000 27920
rect 28533 27915 28599 27918
rect 29200 27888 30000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 841 24714 907 24717
rect 798 24712 907 24714
rect 798 24656 846 24712
rect 902 24656 907 24712
rect 798 24651 907 24656
rect 798 24608 858 24651
rect 0 24518 858 24608
rect 0 24488 800 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 28441 23218 28507 23221
rect 29200 23218 30000 23248
rect 28441 23216 30000 23218
rect 28441 23160 28446 23216
rect 28502 23160 30000 23216
rect 28441 23158 30000 23160
rect 28441 23155 28507 23158
rect 29200 23128 30000 23158
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 28533 22538 28599 22541
rect 29200 22538 30000 22568
rect 28533 22536 30000 22538
rect 28533 22480 28538 22536
rect 28594 22480 30000 22536
rect 28533 22478 30000 22480
rect 28533 22475 28599 22478
rect 29200 22448 30000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 28533 19818 28599 19821
rect 29200 19818 30000 19848
rect 28533 19816 30000 19818
rect 28533 19760 28538 19816
rect 28594 19760 30000 19816
rect 28533 19758 30000 19760
rect 28533 19755 28599 19758
rect 29200 19728 30000 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 28441 16418 28507 16421
rect 29200 16418 30000 16448
rect 28441 16416 30000 16418
rect 28441 16360 28446 16416
rect 28502 16360 30000 16416
rect 28441 16358 30000 16360
rect 28441 16355 28507 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 29200 16328 30000 16358
rect 4870 16287 5186 16288
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 28165 15738 28231 15741
rect 29200 15738 30000 15768
rect 28165 15736 30000 15738
rect 28165 15680 28170 15736
rect 28226 15680 30000 15736
rect 28165 15678 30000 15680
rect 0 15648 800 15678
rect 28165 15675 28231 15678
rect 29200 15648 30000 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 933 9618 999 9621
rect 0 9616 999 9618
rect 0 9560 938 9616
rect 994 9560 999 9616
rect 0 9558 999 9560
rect 0 9528 800 9558
rect 933 9555 999 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 28533 8258 28599 8261
rect 29200 8258 30000 8288
rect 28533 8256 30000 8258
rect 28533 8200 28538 8256
rect 28594 8200 30000 8256
rect 28533 8198 30000 8200
rect 28533 8195 28599 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 29200 8168 30000 8198
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 46816 5188 47376
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1
transform -1 0 25760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1
transform 1 0 25944 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1
transform 1 0 23276 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1
transform 1 0 20056 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1
transform 1 0 18768 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1
transform -1 0 15824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1
transform 1 0 16192 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1
transform -1 0 26864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1
transform -1 0 26220 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1
transform 1 0 24380 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1
transform 1 0 21620 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1
transform -1 0 20608 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1
transform 1 0 18216 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1
transform 1 0 18216 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1
transform 1 0 17480 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1
transform 1 0 14628 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1
transform 1 0 15088 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1
transform 1 0 13892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1
transform 1 0 14628 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1
transform -1 0 14720 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _382_
timestamp 1
transform -1 0 9660 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _383_
timestamp 1
transform 1 0 6808 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _384_
timestamp 1
transform -1 0 10764 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _385_
timestamp 1
transform 1 0 7176 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _386_
timestamp 1
transform 1 0 7176 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _387_
timestamp 1
transform -1 0 6808 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _388_
timestamp 1
transform -1 0 9660 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _389_
timestamp 1
transform 1 0 10304 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _390_
timestamp 1
transform -1 0 9568 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _391_
timestamp 1
transform 1 0 2852 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _392_
timestamp 1
transform -1 0 5888 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _393_
timestamp 1
transform 1 0 5244 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _394_
timestamp 1
transform 1 0 8372 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _395_
timestamp 1
transform 1 0 8280 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _396_
timestamp 1
transform -1 0 9108 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _397_
timestamp 1
transform 1 0 7268 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _398_
timestamp 1
transform -1 0 7268 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _399_
timestamp 1
transform -1 0 6164 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _400_
timestamp 1
transform 1 0 7084 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _401_
timestamp 1
transform -1 0 6992 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _402_
timestamp 1
transform -1 0 7084 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _403_
timestamp 1
transform -1 0 7636 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _404_
timestamp 1
transform 1 0 6716 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _405_
timestamp 1
transform 1 0 2484 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _406_
timestamp 1
transform 1 0 4416 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _407_
timestamp 1
transform -1 0 8280 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _408_
timestamp 1
transform -1 0 6164 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _409_
timestamp 1
transform -1 0 6808 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _410_
timestamp 1
transform -1 0 13616 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _411_
timestamp 1
transform 1 0 11960 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _412_
timestamp 1
transform 1 0 12696 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _413_
timestamp 1
transform 1 0 12512 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _414_
timestamp 1
transform -1 0 13984 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _415_
timestamp 1
transform 1 0 11960 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _416_
timestamp 1
transform -1 0 11960 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _417_
timestamp 1
transform 1 0 8648 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _418_
timestamp 1
transform -1 0 13064 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _419_
timestamp 1
transform 1 0 6900 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _420_
timestamp 1
transform 1 0 8188 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _421_
timestamp 1
transform -1 0 11960 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _422_
timestamp 1
transform -1 0 13524 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _423_
timestamp 1
transform -1 0 15364 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _424_
timestamp 1
transform -1 0 12696 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _425_
timestamp 1
transform 1 0 8372 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _426_
timestamp 1
transform -1 0 8464 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _427_
timestamp 1
transform 1 0 8832 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _428_
timestamp 1
transform 1 0 9476 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _429_
timestamp 1
transform -1 0 10304 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _430_
timestamp 1
transform 1 0 8924 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _431_
timestamp 1
transform 1 0 10120 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _432_
timestamp 1
transform 1 0 10304 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _433_
timestamp 1
transform 1 0 3312 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _434_
timestamp 1
transform 1 0 6348 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _435_
timestamp 1
transform -1 0 12328 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _436_
timestamp 1
transform -1 0 8556 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _437_
timestamp 1
transform 1 0 9476 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _438_
timestamp 1
transform -1 0 13064 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _439_
timestamp 1
transform 1 0 9476 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _440_
timestamp 1
transform -1 0 11408 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _441_
timestamp 1
transform 1 0 9936 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _442_
timestamp 1
transform -1 0 9844 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _443_
timestamp 1
transform -1 0 11408 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _444_
timestamp 1
transform 1 0 10488 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _445_
timestamp 1
transform -1 0 10672 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _446_
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _447_
timestamp 1
transform 1 0 5244 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _448_
timestamp 1
transform -1 0 7728 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _449_
timestamp 1
transform -1 0 10028 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _450_
timestamp 1
transform -1 0 11224 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _451_
timestamp 1
transform 1 0 11776 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _452_
timestamp 1
transform -1 0 12604 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _453_
timestamp 1
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _454_
timestamp 1
transform -1 0 11960 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _455_
timestamp 1
transform 1 0 6256 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _456_
timestamp 1
transform -1 0 10396 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _457_
timestamp 1
transform 1 0 10028 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _458_
timestamp 1
transform 1 0 9292 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _459_
timestamp 1
transform 1 0 10488 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _460_
timestamp 1
transform 1 0 10856 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _461_
timestamp 1
transform 1 0 16928 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _462_
timestamp 1
transform -1 0 19228 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _463_
timestamp 1
transform 1 0 17756 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _464_
timestamp 1
transform -1 0 18492 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _465_
timestamp 1
transform 1 0 18492 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _466_
timestamp 1
transform -1 0 18860 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _467_
timestamp 1
transform -1 0 21436 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _468_
timestamp 1
transform -1 0 20424 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _469_
timestamp 1
transform 1 0 19596 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _470_
timestamp 1
transform 1 0 21068 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _471_
timestamp 1
transform 1 0 21436 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _472_
timestamp 1
transform 1 0 20516 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _473_
timestamp 1
transform 1 0 22816 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _474_
timestamp 1
transform -1 0 23184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _475_
timestamp 1
transform 1 0 22356 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _476_
timestamp 1
transform -1 0 24288 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _477_
timestamp 1
transform -1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _478_
timestamp 1
transform -1 0 23736 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _479_
timestamp 1
transform 1 0 25392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _480_
timestamp 1
transform 1 0 25116 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _481_
timestamp 1
transform 1 0 3036 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _482_
timestamp 1
transform 1 0 5796 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _483_
timestamp 1
transform -1 0 8096 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _484_
timestamp 1
transform -1 0 10120 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _485_
timestamp 1
transform 1 0 8648 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _486_
timestamp 1
transform 1 0 9568 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _487_
timestamp 1
transform 1 0 10212 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _488_
timestamp 1
transform 1 0 10396 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _489_
timestamp 1
transform -1 0 11500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _490_
timestamp 1
transform -1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _491_
timestamp 1
transform -1 0 14628 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _492_
timestamp 1
transform 1 0 10396 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _493_
timestamp 1
transform -1 0 10396 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _494_
timestamp 1
transform 1 0 11684 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _495_
timestamp 1
transform -1 0 12236 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _496_
timestamp 1
transform 1 0 12788 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _497_
timestamp 1
transform -1 0 12696 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _498_
timestamp 1
transform 1 0 11868 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _499_
timestamp 1
transform 1 0 12788 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _500_
timestamp 1
transform 1 0 12512 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _501_
timestamp 1
transform 1 0 12236 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _502_
timestamp 1
transform -1 0 13892 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _503_
timestamp 1
transform 1 0 11776 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _504_
timestamp 1
transform -1 0 12512 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _505_
timestamp 1
transform 1 0 13616 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _506_
timestamp 1
transform 1 0 12236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _507_
timestamp 1
transform -1 0 13064 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _508_
timestamp 1
transform 1 0 12512 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _509_
timestamp 1
transform 1 0 12972 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _510_
timestamp 1
transform 1 0 13432 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _511_
timestamp 1
transform -1 0 14536 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _512_
timestamp 1
transform -1 0 11960 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _513_
timestamp 1
transform 1 0 13524 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _514_
timestamp 1
transform -1 0 14536 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _515_
timestamp 1
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _516_
timestamp 1
transform 1 0 13156 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _517_
timestamp 1
transform -1 0 12972 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _518_
timestamp 1
transform 1 0 13156 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _519_
timestamp 1
transform -1 0 12696 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _520_
timestamp 1
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _521_
timestamp 1
transform -1 0 13524 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _522_
timestamp 1
transform -1 0 13800 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _523_
timestamp 1
transform -1 0 14628 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _524_
timestamp 1
transform -1 0 12512 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _525_
timestamp 1
transform 1 0 12512 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _526_
timestamp 1
transform 1 0 14904 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _527_
timestamp 1
transform 1 0 15548 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _528_
timestamp 1
transform -1 0 16560 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _529_
timestamp 1
transform 1 0 13524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _530_
timestamp 1
transform -1 0 13524 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _531_
timestamp 1
transform 1 0 15364 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _532_
timestamp 1
transform 1 0 16652 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _533_
timestamp 1
transform -1 0 16284 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _534_
timestamp 1
transform -1 0 15824 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _535_
timestamp 1
transform 1 0 15088 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _536_
timestamp 1
transform 1 0 15364 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _537_
timestamp 1
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _538_
timestamp 1
transform 1 0 15732 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _539_
timestamp 1
transform 1 0 13340 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _540_
timestamp 1
transform 1 0 14904 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _541_
timestamp 1
transform 1 0 14536 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _542_
timestamp 1
transform -1 0 15732 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _543_
timestamp 1
transform 1 0 17204 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _544_
timestamp 1
transform 1 0 16652 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_1  _545_
timestamp 1
transform 1 0 13984 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _546_
timestamp 1
transform 1 0 14168 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _547_
timestamp 1
transform 1 0 16008 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _548_
timestamp 1
transform -1 0 18584 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _549_
timestamp 1
transform -1 0 18216 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _550_
timestamp 1
transform -1 0 17388 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _551_
timestamp 1
transform -1 0 16836 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _552_
timestamp 1
transform 1 0 16652 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _553_
timestamp 1
transform 1 0 16836 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _554_
timestamp 1
transform -1 0 16560 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _555_
timestamp 1
transform 1 0 18584 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _556_
timestamp 1
transform 1 0 19596 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _557_
timestamp 1
transform 1 0 19872 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _558_
timestamp 1
transform -1 0 20056 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _559_
timestamp 1
transform -1 0 19872 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _560_
timestamp 1
transform 1 0 20516 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _561_
timestamp 1
transform -1 0 19596 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _562_
timestamp 1
transform 1 0 20976 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _563_
timestamp 1
transform -1 0 21620 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _564_
timestamp 1
transform -1 0 21252 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _565_
timestamp 1
transform 1 0 20424 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _566_
timestamp 1
transform 1 0 20608 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _567_
timestamp 1
transform -1 0 20608 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _568_
timestamp 1
transform -1 0 24288 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _569_
timestamp 1
transform 1 0 23552 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _570_
timestamp 1
transform -1 0 24840 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _571_
timestamp 1
transform 1 0 20424 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _572_
timestamp 1
transform -1 0 20976 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _573_
timestamp 1
transform 1 0 23000 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _574_
timestamp 1
transform 1 0 23276 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _575_
timestamp 1
transform -1 0 23368 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _576_
timestamp 1
transform -1 0 23920 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _577_
timestamp 1
transform -1 0 23736 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _578_
timestamp 1
transform 1 0 22632 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _579_
timestamp 1
transform 1 0 23736 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _580_
timestamp 1
transform -1 0 23644 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _581_
timestamp 1
transform 1 0 26220 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _582_
timestamp 1
transform 1 0 27508 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _583_
timestamp 1
transform -1 0 27508 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _584_
timestamp 1
transform -1 0 24932 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _585_
timestamp 1
transform 1 0 23736 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _586_
timestamp 1
transform 1 0 26220 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _587_
timestamp 1
transform 1 0 26680 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _588_
timestamp 1
transform -1 0 26864 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _589_
timestamp 1
transform 1 0 27508 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _590_
timestamp 1
transform -1 0 27600 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _591_
timestamp 1
transform -1 0 27324 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _592_
timestamp 1
transform 1 0 27140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _593_
timestamp 1
transform -1 0 27140 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _594_
timestamp 1
transform 1 0 13248 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _595_
timestamp 1
transform 1 0 13892 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _596_
timestamp 1
transform -1 0 14996 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _597_
timestamp 1
transform 1 0 14352 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _598_
timestamp 1
transform 1 0 14996 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _599_
timestamp 1
transform 1 0 14720 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_1  _600_
timestamp 1
transform 1 0 13340 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _601_
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _602_
timestamp 1
transform 1 0 15272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _603_
timestamp 1
transform -1 0 16744 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _604_
timestamp 1
transform -1 0 16100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _605_
timestamp 1
transform -1 0 16560 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _606_
timestamp 1
transform 1 0 15272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _607_
timestamp 1
transform 1 0 14812 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _608_
timestamp 1
transform 1 0 15456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _609_
timestamp 1
transform -1 0 15272 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _610_
timestamp 1
transform -1 0 17296 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _611_
timestamp 1
transform 1 0 17480 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _612_
timestamp 1
transform -1 0 18676 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _613_
timestamp 1
transform 1 0 17756 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _614_
timestamp 1
transform 1 0 17940 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _615_
timestamp 1
transform -1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _616_
timestamp 1
transform -1 0 18860 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _617_
timestamp 1
transform 1 0 18676 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _618_
timestamp 1
transform 1 0 19228 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _619_
timestamp 1
transform 1 0 19228 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _620_
timestamp 1
transform -1 0 18952 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _621_
timestamp 1
transform 1 0 21068 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _622_
timestamp 1
transform -1 0 19504 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _623_
timestamp 1
transform -1 0 19964 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _624_
timestamp 1
transform 1 0 21804 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _625_
timestamp 1
transform 1 0 22172 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _626_
timestamp 1
transform -1 0 22172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _627_
timestamp 1
transform 1 0 21068 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _628_
timestamp 1
transform -1 0 22172 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _629_
timestamp 1
transform 1 0 21344 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _630_
timestamp 1
transform 1 0 21988 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _631_
timestamp 1
transform -1 0 21804 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _632_
timestamp 1
transform 1 0 23828 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _633_
timestamp 1
transform 1 0 25024 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _634_
timestamp 1
transform -1 0 25576 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _635_
timestamp 1
transform 1 0 22816 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _636_
timestamp 1
transform -1 0 22816 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _637_
timestamp 1
transform 1 0 24380 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _638_
timestamp 1
transform 1 0 24564 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _639_
timestamp 1
transform -1 0 24012 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _640_
timestamp 1
transform -1 0 25024 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _641_
timestamp 1
transform 1 0 24564 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _642_
timestamp 1
transform -1 0 25852 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _643_
timestamp 1
transform 1 0 24472 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _644_
timestamp 1
transform -1 0 25392 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _645_
timestamp 1
transform 1 0 18216 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _646_
timestamp 1
transform 1 0 17296 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _647_
timestamp 1
transform -1 0 18400 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _648_
timestamp 1
transform 1 0 16652 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _649_
timestamp 1
transform -1 0 16468 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _650_
timestamp 1
transform -1 0 16284 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _651_
timestamp 1
transform 1 0 15640 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _652_
timestamp 1
transform -1 0 15640 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _653_
timestamp 1
transform 1 0 16652 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _654_
timestamp 1
transform -1 0 17940 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _655_
timestamp 1
transform -1 0 17388 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _656_
timestamp 1
transform 1 0 17572 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _657_
timestamp 1
transform 1 0 17572 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _658_
timestamp 1
transform 1 0 17480 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _659_
timestamp 1
transform -1 0 18676 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _660_
timestamp 1
transform 1 0 24564 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _661_
timestamp 1
transform -1 0 19136 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _662_
timestamp 1
transform -1 0 20056 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _663_
timestamp 1
transform 1 0 21068 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _664_
timestamp 1
transform -1 0 20608 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _665_
timestamp 1
transform 1 0 21988 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _666_
timestamp 1
transform 1 0 23460 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _667_
timestamp 1
transform 1 0 25208 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _668_
timestamp 1
transform 1 0 26956 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_1  _669_
timestamp 1
transform 1 0 26312 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _670_
timestamp 1
transform 1 0 15180 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _671_
timestamp 1
transform 1 0 15824 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _672_
timestamp 1
transform 1 0 15640 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _673_
timestamp 1
transform -1 0 16468 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _674_
timestamp 1
transform 1 0 16652 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _675_
timestamp 1
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _676_
timestamp 1
transform 1 0 18308 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _677_
timestamp 1
transform 1 0 18768 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _678_
timestamp 1
transform -1 0 18216 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _679_
timestamp 1
transform -1 0 19688 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _680_
timestamp 1
transform 1 0 19688 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _681_
timestamp 1
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _682_
timestamp 1
transform 1 0 19320 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _683_
timestamp 1
transform 1 0 19780 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _684_
timestamp 1
transform 1 0 18584 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _685_
timestamp 1
transform 1 0 19780 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _686_
timestamp 1
transform -1 0 20516 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _687_
timestamp 1
transform -1 0 22080 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _688_
timestamp 1
transform -1 0 21252 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _689_
timestamp 1
transform -1 0 22632 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _690_
timestamp 1
transform 1 0 24196 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _691_
timestamp 1
transform 1 0 21436 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _692_
timestamp 1
transform -1 0 17572 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _693_
timestamp 1
transform 1 0 17480 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _694_
timestamp 1
transform 1 0 18308 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _695_
timestamp 1
transform -1 0 19872 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _696_
timestamp 1
transform -1 0 21160 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _697_
timestamp 1
transform 1 0 19872 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _698_
timestamp 1
transform 1 0 21896 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _699_
timestamp 1
transform 1 0 23276 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _700_
timestamp 1
transform -1 0 25300 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _701_
timestamp 1
transform -1 0 25944 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _702_
timestamp 1
transform 1 0 17756 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _703_
timestamp 1
transform 1 0 18032 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _704_
timestamp 1
transform -1 0 18952 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _705_
timestamp 1
transform -1 0 19780 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _706_
timestamp 1
transform 1 0 19412 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _707_
timestamp 1
transform 1 0 20700 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _708_
timestamp 1
transform 1 0 21712 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _709_
timestamp 1
transform 1 0 23276 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _710_
timestamp 1
transform -1 0 21712 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _711_
timestamp 1
transform 1 0 22908 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _712_
timestamp 1
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _713_
timestamp 1
transform 1 0 22172 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _714_
timestamp 1
transform -1 0 24932 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _715_
timestamp 1
transform -1 0 24288 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _716_
timestamp 1
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _717_
timestamp 1
transform 1 0 25024 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _718_
timestamp 1
transform 1 0 25484 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _719_
timestamp 1
transform -1 0 25484 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _720_
timestamp 1
transform -1 0 26956 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _721_
timestamp 1
transform -1 0 27048 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _722_
timestamp 1
transform 1 0 8924 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _723_
timestamp 1
transform 1 0 3864 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _724_
timestamp 1
transform 1 0 4784 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _725_
timestamp 1
transform 1 0 5336 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _726_
timestamp 1
transform 1 0 6348 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _727_
timestamp 1
transform 1 0 7360 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _728_
timestamp 1
transform 1 0 8832 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _729_
timestamp 1
transform -1 0 10304 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _730_
timestamp 1
transform 1 0 8924 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _731_
timestamp 1
transform 1 0 7360 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _732_
timestamp 1
transform 1 0 3128 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _733_
timestamp 1
transform 1 0 4692 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _734_
timestamp 1
transform -1 0 7820 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _735_
timestamp 1
transform -1 0 6900 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _736_
timestamp 1
transform 1 0 5244 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _737_
timestamp 1
transform 1 0 5336 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _738_
timestamp 1
transform 1 0 4784 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _739_
timestamp 1
transform 1 0 5428 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _740_
timestamp 1
transform 1 0 12052 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _741_
timestamp 1
transform 1 0 7360 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _742_
timestamp 1
transform 1 0 9200 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _743_
timestamp 1
transform 1 0 9844 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _744_
timestamp 1
transform 1 0 10212 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _745_
timestamp 1
transform 1 0 11040 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _746_
timestamp 1
transform 1 0 12696 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _747_
timestamp 1
transform 1 0 12512 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _748_
timestamp 1
transform -1 0 14628 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _749_
timestamp 1
transform 1 0 10672 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _750_
timestamp 1
transform 1 0 4784 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _751_
timestamp 1
transform 1 0 6808 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _752_
timestamp 1
transform 1 0 9292 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _753_
timestamp 1
transform -1 0 10764 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _754_
timestamp 1
transform 1 0 7268 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _755_
timestamp 1
transform 1 0 7636 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _756_
timestamp 1
transform 1 0 8924 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _757_
timestamp 1
transform 1 0 9568 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _758_
timestamp 1
transform 1 0 12052 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _759_
timestamp 1
transform 1 0 5796 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _760_
timestamp 1
transform 1 0 7176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _761_
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _762_
timestamp 1
transform 1 0 9108 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _763_
timestamp 1
transform -1 0 12880 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _764_
timestamp 1
transform -1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _765_
timestamp 1
transform 1 0 9292 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _766_
timestamp 1
transform -1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _767_
timestamp 1
transform 1 0 11224 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _768_
timestamp 1
transform 1 0 16560 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _769_
timestamp 1
transform -1 0 18124 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _770_
timestamp 1
transform 1 0 18308 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _771_
timestamp 1
transform 1 0 19504 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _772_
timestamp 1
transform 1 0 20148 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _773_
timestamp 1
transform 1 0 21988 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _774_
timestamp 1
transform 1 0 23460 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _775_
timestamp 1
transform 1 0 24932 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _776_
timestamp 1
transform 1 0 8740 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _777_
timestamp 1
transform 1 0 4140 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _778_
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _779_
timestamp 1
transform 1 0 6716 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _780_
timestamp 1
transform 1 0 7268 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _781_
timestamp 1
transform 1 0 9016 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _782_
timestamp 1
transform -1 0 11408 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _783_
timestamp 1
transform -1 0 10580 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _784_
timestamp 1
transform 1 0 8924 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _785_
timestamp 1
transform -1 0 14812 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _786_
timestamp 1
transform 1 0 12420 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _787_
timestamp 1
transform 1 0 11960 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _788_
timestamp 1
transform 1 0 14352 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _789_
timestamp 1
transform 1 0 11224 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _790_
timestamp 1
transform 1 0 12512 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _791_
timestamp 1
transform -1 0 16560 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _792_
timestamp 1
transform -1 0 17112 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _793_
timestamp 1
transform 1 0 12512 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _794_
timestamp 1
transform 1 0 8924 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _795_
timestamp 1
transform -1 0 17204 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _796_
timestamp 1
transform 1 0 16652 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _797_
timestamp 1
transform 1 0 19044 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _798_
timestamp 1
transform 1 0 19872 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _799_
timestamp 1
transform 1 0 22816 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _800_
timestamp 1
transform 1 0 22816 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _801_
timestamp 1
transform 1 0 26956 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _802_
timestamp 1
transform 1 0 26956 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _803_
timestamp 1
transform 1 0 12328 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _804_
timestamp 1
transform 1 0 12144 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _805_
timestamp 1
transform 1 0 14168 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _806_
timestamp 1
transform 1 0 14444 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _807_
timestamp 1
transform 1 0 16928 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _808_
timestamp 1
transform 1 0 19228 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _809_
timestamp 1
transform 1 0 21804 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _810_
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp 1
transform 1 0 24380 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _812_
timestamp 1
transform 1 0 24748 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp 1
transform 1 0 26956 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _814_
timestamp 1
transform 1 0 12052 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _815_
timestamp 1
transform 1 0 26864 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _816_
timestamp 1
transform 1 0 14628 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _817_
timestamp 1
transform 1 0 15272 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _818_
timestamp 1
transform -1 0 17480 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _819_
timestamp 1
transform -1 0 21160 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _820_
timestamp 1
transform 1 0 18216 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _821_
timestamp 1
transform 1 0 19320 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _822_
timestamp 1
transform -1 0 20884 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _823_
timestamp 1
transform -1 0 21252 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _824_
timestamp 1
transform 1 0 26864 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _825_
timestamp 1
transform 1 0 17756 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _826_
timestamp 1
transform -1 0 20700 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _827_
timestamp 1
transform -1 0 21068 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _828_
timestamp 1
transform 1 0 21804 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _829_
timestamp 1
transform 1 0 21804 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _830_
timestamp 1
transform 1 0 23644 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _831_
timestamp 1
transform 1 0 25116 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _832_
timestamp 1
transform 1 0 26956 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _843_
timestamp 1
transform -1 0 27784 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 18032 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1
transform 1 0 8188 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1
transform -1 0 9568 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1
transform -1 0 18768 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1
transform 1 0 17940 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1
transform 1 0 9292 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1
transform -1 0 12328 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1
transform 1 0 19872 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1
transform 1 0 20424 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp 1
transform 1 0 7728 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload2
timestamp 1
transform 1 0 16928 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload3
timestamp 1
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload4
timestamp 1
transform 1 0 10488 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload5
timestamp 1
transform 1 0 20700 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_6  clkload6
timestamp 1
transform 1 0 20424 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1
transform -1 0 16376 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1
transform 1 0 17848 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 1
transform -1 0 17848 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout16
timestamp 1
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1
transform 1 0 13064 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout18
timestamp 1
transform -1 0 12880 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1
transform -1 0 12052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1
transform -1 0 7636 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 1
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 1
transform 1 0 11132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1
transform 1 0 12144 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout26
timestamp 1
transform 1 0 12512 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout27
timestamp 1
transform -1 0 13156 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout28
timestamp 1
transform -1 0 24564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1
transform -1 0 23644 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1
transform -1 0 25760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1
transform -1 0 20976 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 1
transform 1 0 26956 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1
transform -1 0 25944 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_3
timestamp 1562078211
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_15
timestamp 1562078211
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_29
timestamp 1562078211
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_0_41
timestamp 1
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_48
timestamp 1
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_57
timestamp 1562078211
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_69
timestamp 1562078211
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_85
timestamp 1562078211
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_97
timestamp 1562078211
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_113
timestamp 1562078211
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_125
timestamp 1562078211
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_141
timestamp 1562078211
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_153
timestamp 1562078211
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_169
timestamp 1562078211
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_181
timestamp 1562078211
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_197
timestamp 1562078211
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_209
timestamp 1562078211
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_225
timestamp 1562078211
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_237
timestamp 1562078211
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_253
timestamp 1562078211
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_265
timestamp 1562078211
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_286
timestamp 1562078211
transform 1 0 27416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298
timestamp 1
transform 1 0 28520 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_3
timestamp 1562078211
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_15
timestamp 1562078211
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_27
timestamp 1562078211
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_39
timestamp 1562078211
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_57
timestamp 1562078211
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_69
timestamp 1562078211
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_81
timestamp 1562078211
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_93
timestamp 1562078211
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_109
timestamp 1
transform 1 0 11132 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_113
timestamp 1562078211
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_125
timestamp 1562078211
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_137
timestamp 1562078211
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_149
timestamp 1562078211
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_165
timestamp 1
transform 1 0 16284 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_169
timestamp 1562078211
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_181
timestamp 1562078211
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_193
timestamp 1562078211
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_205
timestamp 1562078211
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_225
timestamp 1562078211
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_237
timestamp 1562078211
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_249
timestamp 1562078211
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_261
timestamp 1562078211
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_277
timestamp 1
transform 1 0 26588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_281
timestamp 1562078211
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_293
timestamp 1
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 1
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_3
timestamp 1562078211
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_15
timestamp 1562078211
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_29
timestamp 1562078211
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_41
timestamp 1562078211
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_53
timestamp 1562078211
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_65
timestamp 1562078211
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 1
transform 1 0 8556 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_85
timestamp 1562078211
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_97
timestamp 1562078211
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_109
timestamp 1562078211
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_121
timestamp 1562078211
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_137
timestamp 1
transform 1 0 13708 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_141
timestamp 1562078211
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_153
timestamp 1562078211
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_165
timestamp 1562078211
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_177
timestamp 1562078211
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_193
timestamp 1
transform 1 0 18860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_197
timestamp 1562078211
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_209
timestamp 1562078211
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_221
timestamp 1562078211
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_233
timestamp 1562078211
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_249
timestamp 1
transform 1 0 24012 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_253
timestamp 1562078211
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_265
timestamp 1562078211
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_277
timestamp 1562078211
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_2_289
timestamp 1
transform 1 0 27692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_3
timestamp 1562078211
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_15
timestamp 1562078211
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_27
timestamp 1562078211
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_39
timestamp 1562078211
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_57
timestamp 1562078211
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_69
timestamp 1562078211
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_81
timestamp 1562078211
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_93
timestamp 1562078211
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1
transform 1 0 11132 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_113
timestamp 1562078211
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_125
timestamp 1562078211
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_137
timestamp 1562078211
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_149
timestamp 1562078211
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1
transform 1 0 16284 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_169
timestamp 1562078211
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_181
timestamp 1562078211
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_193
timestamp 1562078211
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_205
timestamp 1562078211
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_225
timestamp 1562078211
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_237
timestamp 1562078211
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_249
timestamp 1562078211
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_261
timestamp 1562078211
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_277
timestamp 1
transform 1 0 26588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_281
timestamp 1562078211
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_293
timestamp 1
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_297
timestamp 1
transform 1 0 28428 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_3
timestamp 1562078211
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_15
timestamp 1562078211
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_29
timestamp 1562078211
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_41
timestamp 1562078211
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_53
timestamp 1562078211
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_65
timestamp 1562078211
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1
transform 1 0 8556 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_85
timestamp 1562078211
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_97
timestamp 1562078211
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_109
timestamp 1562078211
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_121
timestamp 1562078211
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1
transform 1 0 13708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_141
timestamp 1562078211
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_153
timestamp 1562078211
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_165
timestamp 1562078211
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_177
timestamp 1562078211
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1
transform 1 0 18860 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_197
timestamp 1562078211
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_209
timestamp 1562078211
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_221
timestamp 1562078211
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_233
timestamp 1562078211
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_249
timestamp 1
transform 1 0 24012 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_253
timestamp 1562078211
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_265
timestamp 1562078211
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_277
timestamp 1562078211
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_4_289
timestamp 1
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_3
timestamp 1562078211
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_15
timestamp 1562078211
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_27
timestamp 1562078211
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_39
timestamp 1562078211
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_57
timestamp 1562078211
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_69
timestamp 1562078211
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_81
timestamp 1562078211
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_93
timestamp 1562078211
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1
transform 1 0 11132 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_113
timestamp 1562078211
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_125
timestamp 1562078211
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_137
timestamp 1562078211
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_149
timestamp 1562078211
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1
transform 1 0 16284 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_169
timestamp 1562078211
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_181
timestamp 1562078211
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_193
timestamp 1562078211
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_205
timestamp 1562078211
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1
transform 1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_225
timestamp 1562078211
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_237
timestamp 1562078211
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_249
timestamp 1562078211
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_261
timestamp 1562078211
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_277
timestamp 1
transform 1 0 26588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_281
timestamp 1562078211
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_293
timestamp 1
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_3
timestamp 1562078211
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_15
timestamp 1562078211
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_29
timestamp 1562078211
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_41
timestamp 1562078211
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_53
timestamp 1562078211
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_65
timestamp 1562078211
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_81
timestamp 1
transform 1 0 8556 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_85
timestamp 1562078211
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_97
timestamp 1562078211
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_109
timestamp 1562078211
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_121
timestamp 1562078211
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_137
timestamp 1
transform 1 0 13708 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_141
timestamp 1562078211
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_153
timestamp 1562078211
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_165
timestamp 1562078211
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_177
timestamp 1562078211
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_193
timestamp 1
transform 1 0 18860 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_197
timestamp 1562078211
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_209
timestamp 1562078211
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_221
timestamp 1562078211
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_233
timestamp 1562078211
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_249
timestamp 1
transform 1 0 24012 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_253
timestamp 1562078211
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_265
timestamp 1562078211
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_277
timestamp 1562078211
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_6_289
timestamp 1
transform 1 0 27692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_3
timestamp 1562078211
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_15
timestamp 1562078211
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_27
timestamp 1562078211
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_39
timestamp 1562078211
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_57
timestamp 1562078211
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_69
timestamp 1562078211
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_81
timestamp 1562078211
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_93
timestamp 1562078211
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1
transform 1 0 11132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_113
timestamp 1562078211
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_125
timestamp 1562078211
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_137
timestamp 1562078211
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_149
timestamp 1562078211
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_165
timestamp 1
transform 1 0 16284 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_169
timestamp 1562078211
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_181
timestamp 1562078211
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_193
timestamp 1562078211
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_205
timestamp 1562078211
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_225
timestamp 1562078211
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_237
timestamp 1562078211
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_249
timestamp 1562078211
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_261
timestamp 1562078211
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_277
timestamp 1
transform 1 0 26588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_281
timestamp 1562078211
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_293
timestamp 1
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 1
transform 1 0 28428 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_3
timestamp 1562078211
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_15
timestamp 1562078211
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_29
timestamp 1562078211
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_41
timestamp 1562078211
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_53
timestamp 1562078211
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_65
timestamp 1562078211
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_81
timestamp 1
transform 1 0 8556 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_85
timestamp 1562078211
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_97
timestamp 1562078211
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_109
timestamp 1562078211
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_121
timestamp 1562078211
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1
transform 1 0 13708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_141
timestamp 1562078211
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_153
timestamp 1562078211
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_165
timestamp 1562078211
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_177
timestamp 1562078211
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_193
timestamp 1
transform 1 0 18860 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_197
timestamp 1562078211
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_209
timestamp 1562078211
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_221
timestamp 1562078211
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_233
timestamp 1562078211
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_249
timestamp 1
transform 1 0 24012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_253
timestamp 1562078211
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_265
timestamp 1562078211
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_277
timestamp 1562078211
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_8_289
timestamp 1
transform 1 0 27692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_3
timestamp 1562078211
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_15
timestamp 1562078211
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_27
timestamp 1562078211
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_39
timestamp 1562078211
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_51
timestamp 1
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_57
timestamp 1562078211
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_69
timestamp 1562078211
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_81
timestamp 1562078211
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_93
timestamp 1562078211
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_105
timestamp 1
transform 1 0 10764 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1
transform 1 0 11132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_113
timestamp 1562078211
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_125
timestamp 1562078211
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_137
timestamp 1562078211
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_149
timestamp 1562078211
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_169
timestamp 1562078211
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_181
timestamp 1562078211
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_193
timestamp 1562078211
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_205
timestamp 1562078211
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_217
timestamp 1
transform 1 0 21068 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_225
timestamp 1562078211
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_237
timestamp 1562078211
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_249
timestamp 1562078211
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_261
timestamp 1562078211
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_273
timestamp 1
transform 1 0 26220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_277
timestamp 1
transform 1 0 26588 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_281
timestamp 1562078211
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_293
timestamp 1
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_297
timestamp 1
transform 1 0 28428 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_3
timestamp 1562078211
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_15
timestamp 1562078211
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_29
timestamp 1562078211
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_41
timestamp 1562078211
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_53
timestamp 1562078211
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_65
timestamp 1562078211
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_10_77
timestamp 1
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_81
timestamp 1
transform 1 0 8556 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_101
timestamp 1562078211
transform 1 0 10396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_113
timestamp 1562078211
transform 1 0 11500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_125
timestamp 1562078211
transform 1 0 12604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_137
timestamp 1
transform 1 0 13708 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_141
timestamp 1562078211
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_153
timestamp 1562078211
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_165
timestamp 1562078211
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_177
timestamp 1562078211
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_10_189
timestamp 1
transform 1 0 18492 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_193
timestamp 1
transform 1 0 18860 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_213
timestamp 1562078211
transform 1 0 20700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_225
timestamp 1562078211
transform 1 0 21804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_237
timestamp 1562078211
transform 1 0 22908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_249
timestamp 1
transform 1 0 24012 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_253
timestamp 1562078211
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_265
timestamp 1562078211
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_277
timestamp 1562078211
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_10_289
timestamp 1
transform 1 0 27692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_3
timestamp 1562078211
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_15
timestamp 1562078211
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_27
timestamp 1562078211
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_39
timestamp 1
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_43
timestamp 1
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_11_50
timestamp 1
transform 1 0 5704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_11_57
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_65
timestamp 1
transform 1 0 7084 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_72
timestamp 1562078211
transform 1 0 7728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_84
timestamp 1
transform 1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_88
timestamp 1
transform 1 0 9200 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_119
timestamp 1562078211
transform 1 0 12052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_131
timestamp 1562078211
transform 1 0 13156 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_143
timestamp 1
transform 1 0 14260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_147
timestamp 1
transform 1 0 14628 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_154
timestamp 1562078211
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_171
timestamp 1
transform 1 0 16836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1
transform 1 0 18400 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_190
timestamp 1
transform 1 0 18584 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_194
timestamp 1562078211
transform 1 0 18952 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_206
timestamp 1562078211
transform 1 0 20056 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_218
timestamp 1
transform 1 0 21160 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_241
timestamp 1562078211
transform 1 0 23276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_253
timestamp 1562078211
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_265
timestamp 1562078211
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_277
timestamp 1
transform 1 0 26588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_281
timestamp 1562078211
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_293
timestamp 1
transform 1 0 28060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_295
timestamp 1
transform 1 0 28244 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_3
timestamp 1562078211
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_15
timestamp 1562078211
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_29
timestamp 1562078211
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_12_41
timestamp 1
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_49
timestamp 1
transform 1 0 5612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_67
timestamp 1
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_12_77
timestamp 1
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_81
timestamp 1
transform 1 0 8556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_12_85
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_12_98
timestamp 1
transform 1 0 10120 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_125
timestamp 1562078211
transform 1 0 12604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_137
timestamp 1
transform 1 0 13708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_158
timestamp 1562078211
transform 1 0 15640 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_170
timestamp 1
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_174
timestamp 1
transform 1 0 17112 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_178
timestamp 1562078211
transform 1 0 17480 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_190
timestamp 1
transform 1 0 18584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_209
timestamp 1562078211
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_233
timestamp 1562078211
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_245
timestamp 1
transform 1 0 23644 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_249
timestamp 1
transform 1 0 24012 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_269
timestamp 1562078211
transform 1 0 25852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_281
timestamp 1562078211
transform 1 0 26956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_293
timestamp 1
transform 1 0 28060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_3
timestamp 1562078211
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_15
timestamp 1562078211
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_27
timestamp 1562078211
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_39
timestamp 1562078211
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_57
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_82
timestamp 1
transform 1 0 8648 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_90
timestamp 1
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_103
timestamp 1
transform 1 0 10580 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_129
timestamp 1562078211
transform 1 0 12972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_141
timestamp 1
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_148
timestamp 1
transform 1 0 14720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_150
timestamp 1
transform 1 0 14904 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_155
timestamp 1562078211
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_169
timestamp 1562078211
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_181
timestamp 1
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_185
timestamp 1
transform 1 0 18124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_193
timestamp 1
transform 1 0 18860 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_200
timestamp 1562078211
transform 1 0 19504 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_212
timestamp 1
transform 1 0 20608 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_216
timestamp 1
transform 1 0 20976 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_232
timestamp 1562078211
transform 1 0 22448 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_244
timestamp 1
transform 1 0 23552 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_268
timestamp 1562078211
transform 1 0 25760 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_281
timestamp 1562078211
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_293
timestamp 1
transform 1 0 28060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_6
timestamp 1562078211
transform 1 0 1656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_14_18
timestamp 1
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_29
timestamp 1562078211
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_41
timestamp 1562078211
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_53
timestamp 1562078211
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_65
timestamp 1562078211
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_14_77
timestamp 1
transform 1 0 8188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_81
timestamp 1
transform 1 0 8556 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_85
timestamp 1562078211
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_128
timestamp 1562078211
transform 1 0 12880 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_14_141
timestamp 1
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1
transform 1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_154
timestamp 1562078211
transform 1 0 15272 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_166
timestamp 1562078211
transform 1 0 16376 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_204
timestamp 1562078211
transform 1 0 19872 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_216
timestamp 1562078211
transform 1 0 20976 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_228
timestamp 1562078211
transform 1 0 22080 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_14_240
timestamp 1
transform 1 0 23184 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_244
timestamp 1
transform 1 0 23552 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_246
timestamp 1
transform 1 0 23736 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_273
timestamp 1562078211
transform 1 0 26220 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_285
timestamp 1562078211
transform 1 0 27324 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_3
timestamp 1562078211
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_15
timestamp 1562078211
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_27
timestamp 1562078211
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_39
timestamp 1562078211
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_57
timestamp 1562078211
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_69
timestamp 1562078211
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp 1
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_95
timestamp 1562078211
transform 1 0 9844 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_120
timestamp 1
transform 1 0 12144 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_133
timestamp 1562078211
transform 1 0 13340 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_161
timestamp 1
transform 1 0 15916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_165
timestamp 1
transform 1 0 16284 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_169
timestamp 1562078211
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_190
timestamp 1
transform 1 0 18584 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_205
timestamp 1562078211
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_217
timestamp 1
transform 1 0 21068 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_225
timestamp 1562078211
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_237
timestamp 1562078211
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_249
timestamp 1
transform 1 0 24012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_253
timestamp 1
transform 1 0 24380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_265
timestamp 1562078211
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_277
timestamp 1
transform 1 0 26588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_281
timestamp 1562078211
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_293
timestamp 1
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_297
timestamp 1
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_3
timestamp 1562078211
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_15
timestamp 1562078211
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_29
timestamp 1562078211
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_41
timestamp 1562078211
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_53
timestamp 1562078211
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_65
timestamp 1562078211
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_16_77
timestamp 1
transform 1 0 8188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_81
timestamp 1
transform 1 0 8556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_101
timestamp 1
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_107
timestamp 1
transform 1 0 10948 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_116
timestamp 1
transform 1 0 11776 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_118
timestamp 1
transform 1 0 11960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_135
timestamp 1
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_141
timestamp 1
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_170
timestamp 1562078211
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_182
timestamp 1562078211
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_197
timestamp 1562078211
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_209
timestamp 1562078211
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_221
timestamp 1
transform 1 0 21436 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_236
timestamp 1562078211
transform 1 0 22816 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_16_248
timestamp 1
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_253
timestamp 1562078211
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_265
timestamp 1562078211
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_277
timestamp 1562078211
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_16_289
timestamp 1
transform 1 0 27692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_3
timestamp 1562078211
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_15
timestamp 1562078211
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_27
timestamp 1562078211
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_39
timestamp 1562078211
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_17_51
timestamp 1
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_57
timestamp 1562078211
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_69
timestamp 1562078211
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_17_81
timestamp 1
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_85
timestamp 1
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_17_103
timestamp 1
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_121
timestamp 1562078211
transform 1 0 12236 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_133
timestamp 1562078211
transform 1 0 13340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_17_145
timestamp 1
transform 1 0 14444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_153
timestamp 1
transform 1 0 15180 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_17_175
timestamp 1
transform 1 0 17204 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_183
timestamp 1
transform 1 0 17940 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_191
timestamp 1562078211
transform 1 0 18676 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_203
timestamp 1562078211
transform 1 0 19780 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_17_215
timestamp 1
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_225
timestamp 1562078211
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_237
timestamp 1562078211
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_249
timestamp 1562078211
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_261
timestamp 1562078211
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_17_273
timestamp 1
transform 1 0 26220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_277
timestamp 1
transform 1 0 26588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_281
timestamp 1562078211
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_17_293
timestamp 1
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_3
timestamp 1562078211
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_15
timestamp 1562078211
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_29
timestamp 1562078211
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_41
timestamp 1562078211
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_53
timestamp 1562078211
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_65
timestamp 1562078211
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_18_77
timestamp 1
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1
transform 1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_18_85
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_89
timestamp 1
transform 1 0 9292 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_97
timestamp 1562078211
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_109
timestamp 1562078211
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_18_121
timestamp 1
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_18_130
timestamp 1
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_141
timestamp 1562078211
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_18_153
timestamp 1
transform 1 0 15180 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_161
timestamp 1
transform 1 0 15916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1
transform 1 0 16100 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_167
timestamp 1562078211
transform 1 0 16468 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_179
timestamp 1562078211
transform 1 0 17572 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_18_191
timestamp 1
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_197
timestamp 1562078211
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_18_209
timestamp 1
transform 1 0 20332 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_217
timestamp 1
transform 1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1
transform 1 0 21252 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_242
timestamp 1
transform 1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_253
timestamp 1562078211
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_265
timestamp 1562078211
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_277
timestamp 1562078211
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_18_289
timestamp 1
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_3
timestamp 1562078211
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_15
timestamp 1562078211
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_27
timestamp 1562078211
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_39
timestamp 1562078211
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_19_51
timestamp 1
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_57
timestamp 1562078211
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_69
timestamp 1562078211
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_81
timestamp 1562078211
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_93
timestamp 1562078211
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_19_105
timestamp 1
transform 1 0 10764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_109
timestamp 1
transform 1 0 11132 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_113
timestamp 1562078211
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_125
timestamp 1562078211
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_137
timestamp 1562078211
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_149
timestamp 1562078211
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_19_161
timestamp 1
transform 1 0 15916 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_165
timestamp 1
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_176
timestamp 1562078211
transform 1 0 17296 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_188
timestamp 1562078211
transform 1 0 18400 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_200
timestamp 1562078211
transform 1 0 19504 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_19_212
timestamp 1
transform 1 0 20608 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_216
timestamp 1
transform 1 0 20976 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_244
timestamp 1
transform 1 0 23552 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_252
timestamp 1
transform 1 0 24288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_254
timestamp 1
transform 1 0 24472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_269
timestamp 1
transform 1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_277
timestamp 1
transform 1 0 26588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_281
timestamp 1562078211
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_19_293
timestamp 1
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_3
timestamp 1562078211
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_15
timestamp 1562078211
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_29
timestamp 1562078211
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_41
timestamp 1562078211
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_53
timestamp 1562078211
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_65
timestamp 1562078211
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_20_77
timestamp 1
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_81
timestamp 1
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_85
timestamp 1562078211
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_97
timestamp 1562078211
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_109
timestamp 1562078211
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_121
timestamp 1
transform 1 0 12236 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_141
timestamp 1562078211
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_153
timestamp 1
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_20_168
timestamp 1
transform 1 0 16560 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_176
timestamp 1562078211
transform 1 0 17296 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_20_188
timestamp 1
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_197
timestamp 1562078211
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_209
timestamp 1562078211
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_221
timestamp 1
transform 1 0 21436 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_225
timestamp 1562078211
transform 1 0 21804 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_237
timestamp 1562078211
transform 1 0 22908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_249
timestamp 1
transform 1 0 24012 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_281
timestamp 1562078211
transform 1 0 26956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_20_293
timestamp 1
transform 1 0 28060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_3
timestamp 1562078211
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_15
timestamp 1562078211
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_27
timestamp 1562078211
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_39
timestamp 1562078211
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_21_51
timestamp 1
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_57
timestamp 1562078211
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_69
timestamp 1562078211
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_81
timestamp 1562078211
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_93
timestamp 1562078211
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_21_105
timestamp 1
transform 1 0 10764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_109
timestamp 1
transform 1 0 11132 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_113
timestamp 1562078211
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_125
timestamp 1562078211
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_137
timestamp 1562078211
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_149
timestamp 1562078211
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_21_161
timestamp 1
transform 1 0 15916 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_165
timestamp 1
transform 1 0 16284 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_171
timestamp 1
transform 1 0 16836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_192
timestamp 1562078211
transform 1 0 18768 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_204
timestamp 1562078211
transform 1 0 19872 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_21_216
timestamp 1
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_225
timestamp 1562078211
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_237
timestamp 1562078211
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_21_249
timestamp 1
transform 1 0 24012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_257
timestamp 1
transform 1 0 24748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_264
timestamp 1
transform 1 0 25392 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_268
timestamp 1562078211
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_281
timestamp 1562078211
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_21_293
timestamp 1
transform 1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_3
timestamp 1562078211
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_15
timestamp 1562078211
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_29
timestamp 1562078211
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_41
timestamp 1562078211
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_53
timestamp 1562078211
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_22_65
timestamp 1
transform 1 0 7084 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_69
timestamp 1
transform 1 0 7452 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_98
timestamp 1562078211
transform 1 0 10120 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_110
timestamp 1562078211
transform 1 0 11224 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_22_122
timestamp 1
transform 1 0 12328 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_130
timestamp 1
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_132
timestamp 1
transform 1 0 13248 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_149
timestamp 1562078211
transform 1 0 14812 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_22_161
timestamp 1
transform 1 0 15916 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_169
timestamp 1
transform 1 0 16652 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_171
timestamp 1
transform 1 0 16836 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_179
timestamp 1
transform 1 0 17572 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_22_204
timestamp 1
transform 1 0 19872 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_218
timestamp 1562078211
transform 1 0 21160 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_230
timestamp 1562078211
transform 1 0 22264 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_22_242
timestamp 1
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_253
timestamp 1562078211
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_265
timestamp 1562078211
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_277
timestamp 1562078211
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_22_289
timestamp 1
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_3
timestamp 1562078211
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_15
timestamp 1562078211
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_27
timestamp 1562078211
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_39
timestamp 1562078211
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_57
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1
transform 1 0 7084 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_83
timestamp 1
transform 1 0 8740 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_85
timestamp 1
transform 1 0 8924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_23_108
timestamp 1
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_113
timestamp 1562078211
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_125
timestamp 1
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_129
timestamp 1
transform 1 0 12972 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_131
timestamp 1
transform 1 0 13156 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_151
timestamp 1562078211
transform 1 0 14996 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_163
timestamp 1
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_169
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_183
timestamp 1562078211
transform 1 0 17940 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_195
timestamp 1562078211
transform 1 0 19044 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_207
timestamp 1562078211
transform 1 0 20148 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_219
timestamp 1
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_225
timestamp 1
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_233
timestamp 1562078211
transform 1 0 22540 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_245
timestamp 1562078211
transform 1 0 23644 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_257
timestamp 1562078211
transform 1 0 24748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_23_269
timestamp 1
transform 1 0 25852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_277
timestamp 1
transform 1 0 26588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_281
timestamp 1562078211
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_293
timestamp 1
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1
transform 1 0 28428 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_3
timestamp 1562078211
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_24_15
timestamp 1
transform 1 0 2484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1
transform 1 0 2852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_29
timestamp 1562078211
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_41
timestamp 1562078211
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_53
timestamp 1
transform 1 0 5980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_55
timestamp 1
transform 1 0 6164 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_77
timestamp 1
transform 1 0 8188 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_24_96
timestamp 1
transform 1 0 9936 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1
transform 1 0 10304 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_109
timestamp 1
transform 1 0 11132 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_126
timestamp 1562078211
transform 1 0 12696 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_141
timestamp 1562078211
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_153
timestamp 1562078211
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_24_165
timestamp 1
transform 1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_187
timestamp 1
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_24_197
timestamp 1
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_201
timestamp 1
transform 1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_203
timestamp 1
transform 1 0 19780 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_212
timestamp 1
transform 1 0 20608 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_220
timestamp 1
transform 1 0 21344 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_226
timestamp 1562078211
transform 1 0 21896 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_238
timestamp 1562078211
transform 1 0 23000 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_253
timestamp 1562078211
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_265
timestamp 1562078211
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_277
timestamp 1562078211
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_24_289
timestamp 1
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_6
timestamp 1562078211
transform 1 0 1656 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_18
timestamp 1562078211
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_30
timestamp 1
transform 1 0 3864 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_32
timestamp 1
transform 1 0 4048 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_49
timestamp 1
transform 1 0 5612 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_25_73
timestamp 1
transform 1 0 7820 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_113
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_117
timestamp 1
transform 1 0 11868 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_135
timestamp 1562078211
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_147
timestamp 1562078211
transform 1 0 14628 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_25_159
timestamp 1
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_197
timestamp 1562078211
transform 1 0 19228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_209
timestamp 1562078211
transform 1 0 20332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_225
timestamp 1562078211
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_25_237
timestamp 1
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_250
timestamp 1
transform 1 0 24104 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_263
timestamp 1562078211
transform 1 0 25300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_25_275
timestamp 1
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_281
timestamp 1
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_289
timestamp 1
transform 1 0 27692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_291
timestamp 1
transform 1 0 27876 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_3
timestamp 1562078211
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_15
timestamp 1562078211
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_29
timestamp 1562078211
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_26_41
timestamp 1
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_49
timestamp 1
transform 1 0 5612 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_26_58
timestamp 1
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_64
timestamp 1
transform 1 0 6992 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_73
timestamp 1
transform 1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_81
timestamp 1
transform 1 0 8556 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_26_85
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1
transform 1 0 10028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_125
timestamp 1562078211
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_137
timestamp 1
transform 1 0 13708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_141
timestamp 1562078211
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_153
timestamp 1562078211
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_165
timestamp 1
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_167
timestamp 1
transform 1 0 16468 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_184
timestamp 1
transform 1 0 18032 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_197
timestamp 1562078211
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_209
timestamp 1562078211
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_221
timestamp 1562078211
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_233
timestamp 1562078211
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_26_245
timestamp 1
transform 1 0 23644 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_249
timestamp 1
transform 1 0 24012 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_253
timestamp 1
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_261
timestamp 1
transform 1 0 25116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_263
timestamp 1
transform 1 0 25300 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_270
timestamp 1
transform 1 0 25944 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_296
timestamp 1
transform 1 0 28336 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_298
timestamp 1
transform 1 0 28520 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_3
timestamp 1562078211
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_15
timestamp 1562078211
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_27
timestamp 1562078211
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_39
timestamp 1562078211
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_27_51
timestamp 1
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_57
timestamp 1562078211
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_69
timestamp 1562078211
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_81
timestamp 1562078211
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_93
timestamp 1
transform 1 0 9660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_95
timestamp 1
transform 1 0 9844 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_113
timestamp 1562078211
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_125
timestamp 1562078211
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_137
timestamp 1562078211
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_149
timestamp 1562078211
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_27_161
timestamp 1
transform 1 0 15916 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_165
timestamp 1
transform 1 0 16284 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_171
timestamp 1
transform 1 0 16836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_27_175
timestamp 1
transform 1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_225
timestamp 1562078211
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_246
timestamp 1562078211
transform 1 0 23736 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_27_258
timestamp 1
transform 1 0 24840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_262
timestamp 1
transform 1 0 25208 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_268
timestamp 1562078211
transform 1 0 25760 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_281
timestamp 1562078211
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_27_293
timestamp 1
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_3
timestamp 1562078211
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_15
timestamp 1562078211
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_29
timestamp 1562078211
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_41
timestamp 1562078211
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_53
timestamp 1562078211
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_65
timestamp 1562078211
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_28_77
timestamp 1
transform 1 0 8188 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_81
timestamp 1
transform 1 0 8556 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_85
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_95
timestamp 1
transform 1 0 9844 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_101
timestamp 1562078211
transform 1 0 10396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_113
timestamp 1562078211
transform 1 0 11500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_125
timestamp 1562078211
transform 1 0 12604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_137
timestamp 1
transform 1 0 13708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_141
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1
transform 1 0 14444 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_163
timestamp 1562078211
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_175
timestamp 1562078211
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_187
timestamp 1
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_193
timestamp 1
transform 1 0 18860 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_197
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_210
timestamp 1
transform 1 0 20424 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_227
timestamp 1
transform 1 0 21988 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_237
timestamp 1
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_267
timestamp 1
transform 1 0 25668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_269
timestamp 1
transform 1 0 25852 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_286
timestamp 1562078211
transform 1 0 27416 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_298
timestamp 1
transform 1 0 28520 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_3
timestamp 1562078211
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_15
timestamp 1562078211
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_27
timestamp 1562078211
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_39
timestamp 1562078211
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_29_51
timestamp 1
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_57
timestamp 1562078211
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_69
timestamp 1562078211
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_81
timestamp 1
transform 1 0 8556 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_103
timestamp 1
transform 1 0 10580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_113
timestamp 1562078211
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_125
timestamp 1562078211
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_137
timestamp 1562078211
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_29_149
timestamp 1
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_156
timestamp 1
transform 1 0 15456 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_158
timestamp 1
transform 1 0 15640 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_169
timestamp 1562078211
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_29_203
timestamp 1
transform 1 0 19780 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_29_275
timestamp 1
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_281
timestamp 1562078211
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_29_293
timestamp 1
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_297
timestamp 1
transform 1 0 28428 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_3
timestamp 1562078211
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_15
timestamp 1562078211
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_29
timestamp 1562078211
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_30_41
timestamp 1
transform 1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_45
timestamp 1
transform 1 0 5244 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_62
timestamp 1562078211
transform 1 0 6808 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_30_74
timestamp 1
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_101
timestamp 1562078211
transform 1 0 10396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_113
timestamp 1562078211
transform 1 0 11500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_125
timestamp 1562078211
transform 1 0 12604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_137
timestamp 1
transform 1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_141
timestamp 1562078211
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_153
timestamp 1562078211
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_165
timestamp 1562078211
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_177
timestamp 1562078211
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_30_189
timestamp 1
transform 1 0 18492 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_193
timestamp 1
transform 1 0 18860 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_199
timestamp 1
transform 1 0 19412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_224
timestamp 1562078211
transform 1 0 21712 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_245
timestamp 1
transform 1 0 23644 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_249
timestamp 1
transform 1 0 24012 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_253
timestamp 1562078211
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_265
timestamp 1562078211
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_277
timestamp 1562078211
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_30_289
timestamp 1
transform 1 0 27692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_3
timestamp 1562078211
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_15
timestamp 1562078211
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_27
timestamp 1562078211
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_39
timestamp 1
transform 1 0 4692 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_71
timestamp 1562078211
transform 1 0 7636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_83
timestamp 1
transform 1 0 8740 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_93
timestamp 1562078211
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_31_105
timestamp 1
transform 1 0 10764 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_113
timestamp 1562078211
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_125
timestamp 1562078211
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_137
timestamp 1562078211
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_31_149
timestamp 1
transform 1 0 14812 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_157
timestamp 1
transform 1 0 15548 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_31_164
timestamp 1
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_169
timestamp 1562078211
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_181
timestamp 1562078211
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_193
timestamp 1562078211
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_205
timestamp 1562078211
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_31_217
timestamp 1
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_225
timestamp 1562078211
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_237
timestamp 1562078211
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_249
timestamp 1562078211
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_261
timestamp 1562078211
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_31_273
timestamp 1
transform 1 0 26220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_277
timestamp 1
transform 1 0 26588 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_281
timestamp 1562078211
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_31_293
timestamp 1
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1
transform 1 0 28428 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_3
timestamp 1562078211
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_15
timestamp 1562078211
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_29
timestamp 1562078211
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_32_41
timestamp 1
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_45
timestamp 1
transform 1 0 5244 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_71
timestamp 1562078211
transform 1 0 7636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_85
timestamp 1562078211
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_97
timestamp 1562078211
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_109
timestamp 1562078211
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 1
transform 1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_147
timestamp 1
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1
transform 1 0 14996 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_153
timestamp 1
transform 1 0 15180 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_178
timestamp 1562078211
transform 1 0 17480 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_32_190
timestamp 1
transform 1 0 18584 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_197
timestamp 1562078211
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_209
timestamp 1562078211
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_221
timestamp 1562078211
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_233
timestamp 1562078211
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_32_245
timestamp 1
transform 1 0 23644 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_249
timestamp 1
transform 1 0 24012 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_253
timestamp 1562078211
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_265
timestamp 1562078211
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_277
timestamp 1562078211
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_32_289
timestamp 1
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_293
timestamp 1
transform 1 0 28060 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_295
timestamp 1
transform 1 0 28244 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_3
timestamp 1562078211
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_15
timestamp 1562078211
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_27
timestamp 1562078211
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_33_39
timestamp 1
transform 1 0 4692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_47
timestamp 1
transform 1 0 5428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_49
timestamp 1
transform 1 0 5612 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_57
timestamp 1562078211
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_71
timestamp 1
transform 1 0 7636 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_92
timestamp 1562078211
transform 1 0 9568 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_33_104
timestamp 1
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_113
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_132
timestamp 1
transform 1 0 13248 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_33_153
timestamp 1
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_159
timestamp 1
transform 1 0 15732 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_33_164
timestamp 1
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_169
timestamp 1562078211
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_181
timestamp 1562078211
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_193
timestamp 1562078211
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_205
timestamp 1562078211
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_33_217
timestamp 1
transform 1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_225
timestamp 1562078211
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_237
timestamp 1562078211
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_249
timestamp 1562078211
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_261
timestamp 1562078211
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_33_273
timestamp 1
transform 1 0 26220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_277
timestamp 1
transform 1 0 26588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_281
timestamp 1562078211
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_33_293
timestamp 1
transform 1 0 28060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1
transform 1 0 28428 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_3
timestamp 1562078211
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_15
timestamp 1562078211
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_29
timestamp 1562078211
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_41
timestamp 1562078211
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_34_53
timestamp 1
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_61
timestamp 1
transform 1 0 6716 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_71
timestamp 1
transform 1 0 7636 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_34_78
timestamp 1
transform 1 0 8280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_85
timestamp 1562078211
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_97
timestamp 1562078211
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_109
timestamp 1562078211
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_34_121
timestamp 1
transform 1 0 12236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_125
timestamp 1
transform 1 0 12604 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_34_130
timestamp 1
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_141
timestamp 1562078211
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_153
timestamp 1562078211
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_165
timestamp 1562078211
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_177
timestamp 1562078211
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_34_189
timestamp 1
transform 1 0 18492 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_193
timestamp 1
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_197
timestamp 1562078211
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_209
timestamp 1562078211
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_221
timestamp 1562078211
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_233
timestamp 1562078211
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_34_245
timestamp 1
transform 1 0 23644 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_249
timestamp 1
transform 1 0 24012 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_253
timestamp 1562078211
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_265
timestamp 1562078211
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_277
timestamp 1562078211
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_34_289
timestamp 1
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_3
timestamp 1562078211
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_15
timestamp 1562078211
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_27
timestamp 1562078211
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_39
timestamp 1562078211
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_51
timestamp 1
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_57
timestamp 1562078211
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_69
timestamp 1562078211
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_81
timestamp 1562078211
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_93
timestamp 1562078211
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_105
timestamp 1
transform 1 0 10764 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_109
timestamp 1
transform 1 0 11132 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_35_113
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_117
timestamp 1
transform 1 0 11868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_126
timestamp 1562078211
transform 1 0 12696 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_138
timestamp 1562078211
transform 1 0 13800 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_150
timestamp 1562078211
transform 1 0 14904 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_162
timestamp 1
transform 1 0 16008 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_169
timestamp 1562078211
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_181
timestamp 1562078211
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_193
timestamp 1562078211
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_205
timestamp 1562078211
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_217
timestamp 1
transform 1 0 21068 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_221
timestamp 1
transform 1 0 21436 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_225
timestamp 1562078211
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_237
timestamp 1562078211
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_249
timestamp 1562078211
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_261
timestamp 1562078211
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_273
timestamp 1
transform 1 0 26220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_277
timestamp 1
transform 1 0 26588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_281
timestamp 1562078211
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_293
timestamp 1
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_297
timestamp 1
transform 1 0 28428 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_3
timestamp 1562078211
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_15
timestamp 1562078211
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_29
timestamp 1562078211
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_41
timestamp 1562078211
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_36_53
timestamp 1
transform 1 0 5980 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_71
timestamp 1562078211
transform 1 0 7636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_85
timestamp 1562078211
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_97
timestamp 1562078211
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_36_109
timestamp 1
transform 1 0 11132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_113
timestamp 1
transform 1 0 11500 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_36_132
timestamp 1
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_141
timestamp 1562078211
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_36_153
timestamp 1
transform 1 0 15180 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_161
timestamp 1
transform 1 0 15916 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_178
timestamp 1
transform 1 0 17480 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_186
timestamp 1
transform 1 0 18216 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_197
timestamp 1562078211
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_209
timestamp 1562078211
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_221
timestamp 1562078211
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_233
timestamp 1562078211
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_36_245
timestamp 1
transform 1 0 23644 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_249
timestamp 1
transform 1 0 24012 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_253
timestamp 1562078211
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_265
timestamp 1562078211
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_277
timestamp 1562078211
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_36_289
timestamp 1
transform 1 0 27692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_3
timestamp 1562078211
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_15
timestamp 1562078211
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_27
timestamp 1562078211
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_39
timestamp 1562078211
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_37_51
timestamp 1
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_64
timestamp 1
transform 1 0 6992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_68
timestamp 1
transform 1 0 7360 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_77
timestamp 1
transform 1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_81
timestamp 1
transform 1 0 8556 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_87
timestamp 1
transform 1 0 9108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_91
timestamp 1
transform 1 0 9476 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_93
timestamp 1
transform 1 0 9660 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_104
timestamp 1
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_113
timestamp 1562078211
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_125
timestamp 1562078211
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_37_137
timestamp 1
transform 1 0 13708 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_145
timestamp 1
transform 1 0 14444 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_150
timestamp 1562078211
transform 1 0 14904 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_162
timestamp 1
transform 1 0 16008 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp 1
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_179
timestamp 1
transform 1 0 17572 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_218
timestamp 1
transform 1 0 21160 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_225
timestamp 1562078211
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_237
timestamp 1562078211
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_249
timestamp 1562078211
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_261
timestamp 1562078211
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_37_273
timestamp 1
transform 1 0 26220 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_277
timestamp 1
transform 1 0 26588 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_281
timestamp 1562078211
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_293
timestamp 1
transform 1 0 28060 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_295
timestamp 1
transform 1 0 28244 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_3
timestamp 1562078211
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_15
timestamp 1562078211
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_29
timestamp 1562078211
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_38_41
timestamp 1
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_113
timestamp 1
transform 1 0 11500 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_123
timestamp 1562078211
transform 1 0 12420 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_38_135
timestamp 1
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_141
timestamp 1562078211
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_153
timestamp 1562078211
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_38_165
timestamp 1
transform 1 0 16284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_38_178
timestamp 1
transform 1 0 17480 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_186
timestamp 1
transform 1 0 18216 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_188
timestamp 1
transform 1 0 18400 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_213
timestamp 1562078211
transform 1 0 20700 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_225
timestamp 1562078211
transform 1 0 21804 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_237
timestamp 1562078211
transform 1 0 22908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_249
timestamp 1
transform 1 0 24012 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_253
timestamp 1562078211
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_265
timestamp 1562078211
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_38_277
timestamp 1
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_285
timestamp 1
transform 1 0 27324 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_38_290
timestamp 1
transform 1 0 27784 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_298
timestamp 1
transform 1 0 28520 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_3
timestamp 1562078211
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_15
timestamp 1562078211
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_27
timestamp 1562078211
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_39_39
timestamp 1
transform 1 0 4692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_47
timestamp 1
transform 1 0 5428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_49
timestamp 1
transform 1 0 5612 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_70
timestamp 1562078211
transform 1 0 7544 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_39_82
timestamp 1
transform 1 0 8648 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_90
timestamp 1
transform 1 0 9384 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_39_104
timestamp 1
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_113
timestamp 1562078211
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_125
timestamp 1562078211
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_137
timestamp 1562078211
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_149
timestamp 1
transform 1 0 14812 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_176
timestamp 1562078211
transform 1 0 17296 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_39_188
timestamp 1
transform 1 0 18400 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_196
timestamp 1
transform 1 0 19136 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_205
timestamp 1562078211
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_39_217
timestamp 1
transform 1 0 21068 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_221
timestamp 1
transform 1 0 21436 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_225
timestamp 1562078211
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_237
timestamp 1562078211
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_249
timestamp 1562078211
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_261
timestamp 1562078211
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_39_273
timestamp 1
transform 1 0 26220 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_277
timestamp 1
transform 1 0 26588 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_281
timestamp 1562078211
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_293
timestamp 1
transform 1 0 28060 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_3
timestamp 1562078211
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_15
timestamp 1562078211
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_40_29
timestamp 1
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_33
timestamp 1
transform 1 0 4140 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_35
timestamp 1
transform 1 0 4324 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_49
timestamp 1
transform 1 0 5612 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_40_78
timestamp 1
transform 1 0 8280 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_85
timestamp 1562078211
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_97
timestamp 1562078211
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_109
timestamp 1562078211
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_40_121
timestamp 1
transform 1 0 12236 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_129
timestamp 1
transform 1 0 12972 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_131
timestamp 1
transform 1 0 13156 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_141
timestamp 1562078211
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_153
timestamp 1562078211
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_165
timestamp 1562078211
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_177
timestamp 1562078211
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_40_189
timestamp 1
transform 1 0 18492 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_193
timestamp 1
transform 1 0 18860 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_197
timestamp 1562078211
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_209
timestamp 1562078211
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_221
timestamp 1562078211
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_233
timestamp 1562078211
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_40_245
timestamp 1
transform 1 0 23644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_249
timestamp 1
transform 1 0 24012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_253
timestamp 1562078211
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_265
timestamp 1562078211
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_277
timestamp 1562078211
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_40_289
timestamp 1
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_41_6
timestamp 1
transform 1 0 1656 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_14
timestamp 1
transform 1 0 2392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_20
timestamp 1
transform 1 0 2944 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_38
timestamp 1
transform 1 0 4600 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_73
timestamp 1
transform 1 0 7820 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_81
timestamp 1
transform 1 0 8556 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_99
timestamp 1562078211
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_113
timestamp 1562078211
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_41_125
timestamp 1
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_133
timestamp 1
transform 1 0 13340 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_142
timestamp 1562078211
transform 1 0 14168 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_154
timestamp 1562078211
transform 1 0 15272 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_169
timestamp 1562078211
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_181
timestamp 1562078211
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_193
timestamp 1562078211
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_205
timestamp 1562078211
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_41_217
timestamp 1
transform 1 0 21068 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_221
timestamp 1
transform 1 0 21436 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_225
timestamp 1562078211
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_237
timestamp 1562078211
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_249
timestamp 1562078211
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_261
timestamp 1562078211
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_41_273
timestamp 1
transform 1 0 26220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_277
timestamp 1
transform 1 0 26588 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_281
timestamp 1562078211
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_41_293
timestamp 1
transform 1 0 28060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_297
timestamp 1
transform 1 0 28428 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_3
timestamp 1562078211
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_15
timestamp 1562078211
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_29
timestamp 1562078211
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_42_41
timestamp 1
transform 1 0 4876 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_45
timestamp 1
transform 1 0 5244 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_71
timestamp 1562078211
transform 1 0 7636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_85
timestamp 1562078211
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_97
timestamp 1562078211
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_109
timestamp 1562078211
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_42_134
timestamp 1
transform 1 0 13432 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_141
timestamp 1562078211
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_42_153
timestamp 1
transform 1 0 15180 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_161
timestamp 1
transform 1 0 15916 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_165
timestamp 1562078211
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_177
timestamp 1562078211
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_42_189
timestamp 1
transform 1 0 18492 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_193
timestamp 1
transform 1 0 18860 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_197
timestamp 1562078211
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_209
timestamp 1562078211
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_221
timestamp 1562078211
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_233
timestamp 1562078211
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_42_245
timestamp 1
transform 1 0 23644 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_249
timestamp 1
transform 1 0 24012 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_253
timestamp 1562078211
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_265
timestamp 1562078211
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_277
timestamp 1562078211
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_42_289
timestamp 1
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_3
timestamp 1562078211
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_15
timestamp 1562078211
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_27
timestamp 1562078211
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_39
timestamp 1562078211
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_43_51
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_57
timestamp 1562078211
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_69
timestamp 1562078211
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_43_81
timestamp 1
transform 1 0 8556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_85
timestamp 1
transform 1 0 8924 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_87
timestamp 1
transform 1 0 9108 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_93
timestamp 1562078211
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_43_105
timestamp 1
transform 1 0 10764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_109
timestamp 1
transform 1 0 11132 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_115
timestamp 1
transform 1 0 11684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_140
timestamp 1562078211
transform 1 0 13984 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_43_152
timestamp 1
transform 1 0 15088 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_160
timestamp 1
transform 1 0 15824 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_188
timestamp 1562078211
transform 1 0 18400 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_200
timestamp 1562078211
transform 1 0 19504 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_212
timestamp 1562078211
transform 1 0 20608 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_225
timestamp 1562078211
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_237
timestamp 1562078211
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_249
timestamp 1562078211
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_261
timestamp 1562078211
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_43_273
timestamp 1
transform 1 0 26220 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_277
timestamp 1
transform 1 0 26588 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_281
timestamp 1562078211
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_43_293
timestamp 1
transform 1 0 28060 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_297
timestamp 1
transform 1 0 28428 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_3
timestamp 1562078211
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_15
timestamp 1562078211
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_29
timestamp 1562078211
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_41
timestamp 1562078211
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_53
timestamp 1562078211
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_65
timestamp 1562078211
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_44_77
timestamp 1
transform 1 0 8188 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_81
timestamp 1
transform 1 0 8556 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_85
timestamp 1562078211
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_97
timestamp 1562078211
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_44_109
timestamp 1
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_117
timestamp 1
transform 1 0 11868 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_143
timestamp 1
transform 1 0 14260 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_44_160
timestamp 1
transform 1 0 15824 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_184
timestamp 1562078211
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_197
timestamp 1
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_211
timestamp 1562078211
transform 1 0 20516 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_223
timestamp 1562078211
transform 1 0 21620 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_235
timestamp 1562078211
transform 1 0 22724 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_44_247
timestamp 1
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_253
timestamp 1562078211
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_265
timestamp 1562078211
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_277
timestamp 1562078211
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_44_289
timestamp 1
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_3
timestamp 1562078211
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_15
timestamp 1562078211
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_27
timestamp 1562078211
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_39
timestamp 1562078211
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_57
timestamp 1562078211
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_69
timestamp 1562078211
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_45_81
timestamp 1
transform 1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_45_101
timestamp 1
transform 1 0 10396 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_109
timestamp 1
transform 1 0 11132 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_113
timestamp 1
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_121
timestamp 1
transform 1 0 12236 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_123
timestamp 1
transform 1 0 12420 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_146
timestamp 1562078211
transform 1 0 14536 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_45_158
timestamp 1
transform 1 0 15640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_45_169
timestamp 1
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_173
timestamp 1
transform 1 0 17020 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_175
timestamp 1
transform 1 0 17204 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_181
timestamp 1562078211
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_193
timestamp 1
transform 1 0 18860 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_45_219
timestamp 1
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_225
timestamp 1562078211
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_237
timestamp 1562078211
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_249
timestamp 1562078211
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_261
timestamp 1562078211
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_45_273
timestamp 1
transform 1 0 26220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_277
timestamp 1
transform 1 0 26588 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_281
timestamp 1562078211
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_45_293
timestamp 1
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1
transform 1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_3
timestamp 1562078211
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_15
timestamp 1562078211
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_29
timestamp 1562078211
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_41
timestamp 1562078211
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_53
timestamp 1562078211
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_65
timestamp 1562078211
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_46_77
timestamp 1
transform 1 0 8188 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_81
timestamp 1
transform 1 0 8556 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_85
timestamp 1562078211
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_97
timestamp 1562078211
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_109
timestamp 1562078211
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_121
timestamp 1562078211
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_133
timestamp 1
transform 1 0 13340 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_137
timestamp 1
transform 1 0 13708 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_141
timestamp 1562078211
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_153
timestamp 1562078211
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_46_165
timestamp 1
transform 1 0 16284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_175
timestamp 1
transform 1 0 17204 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_186
timestamp 1
transform 1 0 18216 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_197
timestamp 1
transform 1 0 19228 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_234
timestamp 1562078211
transform 1 0 22632 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_46_246
timestamp 1
transform 1 0 23736 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_253
timestamp 1562078211
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_265
timestamp 1562078211
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_277
timestamp 1562078211
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_46_289
timestamp 1
transform 1 0 27692 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_3
timestamp 1562078211
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_15
timestamp 1562078211
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_27
timestamp 1562078211
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_39
timestamp 1562078211
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_57
timestamp 1562078211
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_69
timestamp 1562078211
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_81
timestamp 1562078211
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_93
timestamp 1562078211
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_47_105
timestamp 1
transform 1 0 10764 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_109
timestamp 1
transform 1 0 11132 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_113
timestamp 1562078211
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_125
timestamp 1562078211
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_137
timestamp 1562078211
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_149
timestamp 1562078211
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_47_161
timestamp 1
transform 1 0 15916 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_165
timestamp 1
transform 1 0 16284 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_169
timestamp 1
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_177
timestamp 1
transform 1 0 17388 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_186
timestamp 1562078211
transform 1 0 18216 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_198
timestamp 1
transform 1 0 19320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_225
timestamp 1562078211
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_237
timestamp 1562078211
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_249
timestamp 1562078211
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_261
timestamp 1562078211
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_47_273
timestamp 1
transform 1 0 26220 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_277
timestamp 1
transform 1 0 26588 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_281
timestamp 1562078211
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_293
timestamp 1
transform 1 0 28060 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_295
timestamp 1
transform 1 0 28244 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_3
timestamp 1562078211
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_15
timestamp 1562078211
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_29
timestamp 1562078211
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_41
timestamp 1562078211
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_53
timestamp 1562078211
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_65
timestamp 1562078211
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_48_77
timestamp 1
transform 1 0 8188 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_81
timestamp 1
transform 1 0 8556 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_92
timestamp 1562078211
transform 1 0 9568 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_104
timestamp 1562078211
transform 1 0 10672 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_116
timestamp 1562078211
transform 1 0 11776 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_128
timestamp 1562078211
transform 1 0 12880 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_141
timestamp 1562078211
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_153
timestamp 1562078211
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_165
timestamp 1562078211
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_177
timestamp 1
transform 1 0 17388 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_48_191
timestamp 1
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_48_197
timestamp 1
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_201
timestamp 1
transform 1 0 19596 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_48_206
timestamp 1
transform 1 0 20056 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_214
timestamp 1
transform 1 0 20792 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_219
timestamp 1562078211
transform 1 0 21252 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_231
timestamp 1562078211
transform 1 0 22356 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_48_243
timestamp 1
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_253
timestamp 1562078211
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_265
timestamp 1562078211
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_277
timestamp 1562078211
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_48_289
timestamp 1
transform 1 0 27692 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_297
timestamp 1
transform 1 0 28428 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_6
timestamp 1562078211
transform 1 0 1656 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_18
timestamp 1562078211
transform 1 0 2760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_30
timestamp 1562078211
transform 1 0 3864 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_49_42
timestamp 1
transform 1 0 4968 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_46
timestamp 1
transform 1 0 5336 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_49_57
timestamp 1
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_65
timestamp 1
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_71
timestamp 1
transform 1 0 7636 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_106
timestamp 1
transform 1 0 10856 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_113
timestamp 1562078211
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_125
timestamp 1562078211
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_137
timestamp 1562078211
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_149
timestamp 1
transform 1 0 14812 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_151
timestamp 1
transform 1 0 14996 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_155
timestamp 1562078211
transform 1 0 15364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_169
timestamp 1562078211
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_49_181
timestamp 1
transform 1 0 17756 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_185
timestamp 1
transform 1 0 18124 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_191
timestamp 1562078211
transform 1 0 18676 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_203
timestamp 1562078211
transform 1 0 19780 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_49_215
timestamp 1
transform 1 0 20884 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_225
timestamp 1562078211
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_237
timestamp 1562078211
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_249
timestamp 1562078211
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_261
timestamp 1562078211
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_49_273
timestamp 1
transform 1 0 26220 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_277
timestamp 1
transform 1 0 26588 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_281
timestamp 1562078211
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_49_293
timestamp 1
transform 1 0 28060 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_297
timestamp 1
transform 1 0 28428 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_6
timestamp 1562078211
transform 1 0 1656 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_18
timestamp 1
transform 1 0 2760 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_50_24
timestamp 1
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_29
timestamp 1
transform 1 0 3772 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_113
timestamp 1562078211
transform 1 0 11500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_125
timestamp 1562078211
transform 1 0 12604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_137
timestamp 1
transform 1 0 13708 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_141
timestamp 1562078211
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_50_153
timestamp 1
transform 1 0 15180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_157
timestamp 1
transform 1 0 15548 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_174
timestamp 1562078211
transform 1 0 17112 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_50_186
timestamp 1
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_197
timestamp 1562078211
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_209
timestamp 1562078211
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_221
timestamp 1562078211
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_233
timestamp 1562078211
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_50_245
timestamp 1
transform 1 0 23644 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_249
timestamp 1
transform 1 0 24012 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_253
timestamp 1562078211
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_265
timestamp 1562078211
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_277
timestamp 1562078211
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_50_289
timestamp 1
transform 1 0 27692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_297
timestamp 1
transform 1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_3
timestamp 1562078211
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_15
timestamp 1562078211
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_27
timestamp 1562078211
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_39
timestamp 1
transform 1 0 4692 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_81
timestamp 1
transform 1 0 8556 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_83
timestamp 1
transform 1 0 8740 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_105
timestamp 1
transform 1 0 10764 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_109
timestamp 1
transform 1 0 11132 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_113
timestamp 1562078211
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_125
timestamp 1562078211
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_137
timestamp 1562078211
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_149
timestamp 1
transform 1 0 14812 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_151
timestamp 1
transform 1 0 14996 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_169
timestamp 1562078211
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_181
timestamp 1562078211
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_193
timestamp 1562078211
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_205
timestamp 1562078211
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_51_217
timestamp 1
transform 1 0 21068 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_221
timestamp 1
transform 1 0 21436 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_225
timestamp 1562078211
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_237
timestamp 1562078211
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_249
timestamp 1562078211
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_261
timestamp 1562078211
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_51_273
timestamp 1
transform 1 0 26220 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_277
timestamp 1
transform 1 0 26588 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 1
transform 1 0 28428 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_6
timestamp 1562078211
transform 1 0 1656 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_52_18
timestamp 1
transform 1 0 2760 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_29
timestamp 1562078211
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_52_41
timestamp 1
transform 1 0 4876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_52_73
timestamp 1
transform 1 0 7820 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_81
timestamp 1
transform 1 0 8556 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_85
timestamp 1562078211
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_97
timestamp 1562078211
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_109
timestamp 1
transform 1 0 11132 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_129
timestamp 1
transform 1 0 12972 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_137
timestamp 1
transform 1 0 13708 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_141
timestamp 1562078211
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_153
timestamp 1
transform 1 0 15180 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_162
timestamp 1562078211
transform 1 0 16008 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_174
timestamp 1562078211
transform 1 0 17112 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_52_186
timestamp 1
transform 1 0 18216 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_197
timestamp 1562078211
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_209
timestamp 1562078211
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_221
timestamp 1562078211
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_233
timestamp 1562078211
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_52_245
timestamp 1
transform 1 0 23644 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_249
timestamp 1
transform 1 0 24012 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_253
timestamp 1562078211
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_265
timestamp 1562078211
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_277
timestamp 1562078211
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_52_289
timestamp 1
transform 1 0 27692 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_297
timestamp 1
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_3
timestamp 1562078211
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_15
timestamp 1562078211
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_27
timestamp 1562078211
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_53_39
timestamp 1
transform 1 0 4692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_52
timestamp 1
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_62
timestamp 1562078211
transform 1 0 6808 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_53_74
timestamp 1
transform 1 0 7912 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_91
timestamp 1562078211
transform 1 0 9476 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_53_103
timestamp 1
transform 1 0 10580 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_136
timestamp 1562078211
transform 1 0 13616 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_148
timestamp 1562078211
transform 1 0 14720 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_53_160
timestamp 1
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_169
timestamp 1562078211
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_181
timestamp 1562078211
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_193
timestamp 1562078211
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_205
timestamp 1562078211
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_53_217
timestamp 1
transform 1 0 21068 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_221
timestamp 1
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_225
timestamp 1562078211
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_237
timestamp 1562078211
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_53_249
timestamp 1
transform 1 0 24012 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_257
timestamp 1
transform 1 0 24748 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_268
timestamp 1562078211
transform 1 0 25760 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_281
timestamp 1562078211
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_53_293
timestamp 1
transform 1 0 28060 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 1
transform 1 0 28428 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_6
timestamp 1562078211
transform 1 0 1656 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_54_18
timestamp 1
transform 1 0 2760 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_29
timestamp 1562078211
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_41
timestamp 1562078211
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_53
timestamp 1562078211
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_65
timestamp 1562078211
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_54_77
timestamp 1
transform 1 0 8188 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_81
timestamp 1
transform 1 0 8556 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_101
timestamp 1562078211
transform 1 0 10396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_113
timestamp 1
transform 1 0 11500 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_146
timestamp 1562078211
transform 1 0 14536 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_158
timestamp 1562078211
transform 1 0 15640 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_170
timestamp 1562078211
transform 1 0 16744 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_182
timestamp 1562078211
transform 1 0 17848 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_197
timestamp 1562078211
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_209
timestamp 1562078211
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_221
timestamp 1562078211
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_233
timestamp 1562078211
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_54_245
timestamp 1
transform 1 0 23644 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_267
timestamp 1
transform 1 0 25668 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_282
timestamp 1562078211
transform 1 0 27048 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_294
timestamp 1
transform 1 0 28152 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_6
timestamp 1562078211
transform 1 0 1656 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_18
timestamp 1562078211
transform 1 0 2760 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_30
timestamp 1562078211
transform 1 0 3864 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_42
timestamp 1562078211
transform 1 0 4968 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_57
timestamp 1562078211
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_69
timestamp 1562078211
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_81
timestamp 1562078211
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_93
timestamp 1562078211
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_55_105
timestamp 1
transform 1 0 10764 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_109
timestamp 1
transform 1 0 11132 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_55_113
timestamp 1
transform 1 0 11500 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_117
timestamp 1
transform 1 0 11868 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_126
timestamp 1
transform 1 0 12696 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_150
timestamp 1562078211
transform 1 0 14904 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_55_162
timestamp 1
transform 1 0 16008 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_169
timestamp 1562078211
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_181
timestamp 1562078211
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_55_193
timestamp 1
transform 1 0 18860 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_55_205
timestamp 1
transform 1 0 19964 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_217
timestamp 1
transform 1 0 21068 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_221
timestamp 1
transform 1 0 21436 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_55_225
timestamp 1
transform 1 0 21804 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_55_235
timestamp 1
transform 1 0 22724 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_243
timestamp 1
transform 1 0 23460 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_277
timestamp 1
transform 1 0 26588 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_297
timestamp 1
transform 1 0 28428 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_6
timestamp 1562078211
transform 1 0 1656 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_56_18
timestamp 1
transform 1 0 2760 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_29
timestamp 1562078211
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_41
timestamp 1562078211
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_53
timestamp 1562078211
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_65
timestamp 1562078211
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_56_77
timestamp 1
transform 1 0 8188 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_81
timestamp 1
transform 1 0 8556 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_85
timestamp 1562078211
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_97
timestamp 1562078211
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_109
timestamp 1562078211
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_141
timestamp 1562078211
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_153
timestamp 1
transform 1 0 15180 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_160
timestamp 1562078211
transform 1 0 15824 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_172
timestamp 1562078211
transform 1 0 16928 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_56_184
timestamp 1
transform 1 0 18032 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_56_197
timestamp 1
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_217
timestamp 1
transform 1 0 21068 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_224
timestamp 1
transform 1 0 21712 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_253
timestamp 1
transform 1 0 24380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_259
timestamp 1
transform 1 0 24932 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_265
timestamp 1562078211
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_285
timestamp 1
transform 1 0 27324 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_287
timestamp 1
transform 1 0 27508 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_296
timestamp 1
transform 1 0 28336 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_298
timestamp 1
transform 1 0 28520 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_3
timestamp 1562078211
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_57_15
timestamp 1
transform 1 0 2484 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_23
timestamp 1
transform 1 0 3220 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_29
timestamp 1562078211
transform 1 0 3772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_41
timestamp 1562078211
transform 1 0 4876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_53
timestamp 1
transform 1 0 5980 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_57
timestamp 1562078211
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_69
timestamp 1562078211
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_81
timestamp 1562078211
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_93
timestamp 1562078211
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_57_105
timestamp 1
transform 1 0 10764 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_109
timestamp 1
transform 1 0 11132 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_113
timestamp 1
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_121
timestamp 1
transform 1 0 12236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_123
timestamp 1
transform 1 0 12420 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_148
timestamp 1
transform 1 0 14720 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_197
timestamp 1
transform 1 0 19228 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_244
timestamp 1562078211
transform 1 0 23552 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_256
timestamp 1562078211
transform 1 0 24656 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_268
timestamp 1562078211
transform 1 0 25760 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_281
timestamp 1562078211
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_57_293
timestamp 1
transform 1 0 28060 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_297
timestamp 1
transform 1 0 28428 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_3
timestamp 1562078211
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_15
timestamp 1562078211
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_29
timestamp 1562078211
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_41
timestamp 1562078211
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_53
timestamp 1562078211
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_65
timestamp 1562078211
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_58_77
timestamp 1
transform 1 0 8188 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_81
timestamp 1
transform 1 0 8556 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_85
timestamp 1562078211
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_97
timestamp 1562078211
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_109
timestamp 1562078211
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_121
timestamp 1562078211
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_58_133
timestamp 1
transform 1 0 13340 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_137
timestamp 1
transform 1 0 13708 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_141
timestamp 1562078211
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_58_153
timestamp 1
transform 1 0 15180 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_165
timestamp 1562078211
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_58_177
timestamp 1
transform 1 0 17388 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_58_242
timestamp 1
transform 1 0 23368 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_58_253
timestamp 1
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_261
timestamp 1
transform 1 0 25116 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_269
timestamp 1562078211
transform 1 0 25852 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_58_281
timestamp 1
transform 1 0 26956 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_285
timestamp 1
transform 1 0 27324 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_58_294
timestamp 1
transform 1 0 28152 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_298
timestamp 1
transform 1 0 28520 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_3
timestamp 1562078211
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_15
timestamp 1562078211
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_27
timestamp 1562078211
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_39
timestamp 1
transform 1 0 4692 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_57
timestamp 1562078211
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_69
timestamp 1562078211
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_59_81
timestamp 1
transform 1 0 8556 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_105
timestamp 1
transform 1 0 10764 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_109
timestamp 1
transform 1 0 11132 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_113
timestamp 1562078211
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_125
timestamp 1562078211
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_137
timestamp 1562078211
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_149
timestamp 1
transform 1 0 14812 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_151
timestamp 1
transform 1 0 14996 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_169
timestamp 1562078211
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_59_181
timestamp 1
transform 1 0 17756 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_196
timestamp 1
transform 1 0 19136 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_200
timestamp 1
transform 1 0 19504 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_59_236
timestamp 1
transform 1 0 22816 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_240
timestamp 1
transform 1 0 23184 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_242
timestamp 1
transform 1 0 23368 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_59_251
timestamp 1
transform 1 0 24196 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_260
timestamp 1562078211
transform 1 0 25024 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_272
timestamp 1
transform 1 0 26128 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_59_290
timestamp 1
transform 1 0 27784 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_298
timestamp 1
transform 1 0 28520 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_3
timestamp 1562078211
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_15
timestamp 1562078211
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_29
timestamp 1562078211
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_41
timestamp 1562078211
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_60_53
timestamp 1
transform 1 0 5980 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_65
timestamp 1562078211
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_77
timestamp 1
transform 1 0 8188 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_60_85
timestamp 1
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_122
timestamp 1562078211
transform 1 0 12328 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_60_134
timestamp 1
transform 1 0 13432 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_141
timestamp 1562078211
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_153
timestamp 1562078211
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_165
timestamp 1562078211
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_177
timestamp 1562078211
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_60_189
timestamp 1
transform 1 0 18492 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_193
timestamp 1
transform 1 0 18860 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_216
timestamp 1562078211
transform 1 0 20976 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_228
timestamp 1562078211
transform 1 0 22080 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_240
timestamp 1562078211
transform 1 0 23184 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_253
timestamp 1562078211
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_265
timestamp 1562078211
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_277
timestamp 1
transform 1 0 26588 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_279
timestamp 1
transform 1 0 26772 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_296
timestamp 1
transform 1 0 28336 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_298
timestamp 1
transform 1 0 28520 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_3
timestamp 1562078211
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_15
timestamp 1562078211
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_27
timestamp 1562078211
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_39
timestamp 1562078211
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_61_51
timestamp 1
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_61_78
timestamp 1
transform 1 0 8280 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_82
timestamp 1
transform 1 0 8648 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_61_105
timestamp 1
transform 1 0 10764 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_109
timestamp 1
transform 1 0 11132 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_113
timestamp 1562078211
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_125
timestamp 1562078211
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_137
timestamp 1562078211
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_149
timestamp 1562078211
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_61_161
timestamp 1
transform 1 0 15916 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_165
timestamp 1
transform 1 0 16284 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_169
timestamp 1562078211
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_181
timestamp 1562078211
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_61_193
timestamp 1
transform 1 0 18860 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_197
timestamp 1
transform 1 0 19228 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_203
timestamp 1562078211
transform 1 0 19780 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_61_215
timestamp 1
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_225
timestamp 1562078211
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_237
timestamp 1562078211
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_249
timestamp 1562078211
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_261
timestamp 1562078211
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_61_273
timestamp 1
transform 1 0 26220 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_277
timestamp 1
transform 1 0 26588 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_61_289
timestamp 1
transform 1 0 27692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_293
timestamp 1
transform 1 0 28060 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_3
timestamp 1562078211
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_15
timestamp 1562078211
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_29
timestamp 1562078211
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_41
timestamp 1562078211
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_53
timestamp 1562078211
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_65
timestamp 1562078211
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_62_77
timestamp 1
transform 1 0 8188 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_81
timestamp 1
transform 1 0 8556 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_93
timestamp 1562078211
transform 1 0 9660 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_105
timestamp 1562078211
transform 1 0 10764 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_117
timestamp 1562078211
transform 1 0 11868 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_62_129
timestamp 1
transform 1 0 12972 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_137
timestamp 1
transform 1 0 13708 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_141
timestamp 1562078211
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_153
timestamp 1562078211
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_165
timestamp 1562078211
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_177
timestamp 1562078211
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_62_189
timestamp 1
transform 1 0 18492 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_193
timestamp 1
transform 1 0 18860 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_197
timestamp 1562078211
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_209
timestamp 1
transform 1 0 20332 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_230
timestamp 1562078211
transform 1 0 22264 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_62_242
timestamp 1
transform 1 0 23368 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_253
timestamp 1562078211
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_265
timestamp 1562078211
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_277
timestamp 1562078211
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_62_289
timestamp 1
transform 1 0 27692 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_297
timestamp 1
transform 1 0 28428 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_3
timestamp 1562078211
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_15
timestamp 1562078211
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_27
timestamp 1562078211
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_39
timestamp 1562078211
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_63_51
timestamp 1
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_57
timestamp 1562078211
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_63_69
timestamp 1
transform 1 0 7452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_73
timestamp 1
transform 1 0 7820 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_63_80
timestamp 1
transform 1 0 8464 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_107
timestamp 1
transform 1 0 10948 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_113
timestamp 1
transform 1 0 11500 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_126
timestamp 1562078211
transform 1 0 12696 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_138
timestamp 1562078211
transform 1 0 13800 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_150
timestamp 1562078211
transform 1 0 14904 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_63_162
timestamp 1
transform 1 0 16008 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_169
timestamp 1562078211
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_181
timestamp 1562078211
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_193
timestamp 1562078211
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_63_205
timestamp 1
transform 1 0 19964 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_209
timestamp 1
transform 1 0 20332 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_63_217
timestamp 1
transform 1 0 21068 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_221
timestamp 1
transform 1 0 21436 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_225
timestamp 1562078211
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_237
timestamp 1
transform 1 0 22908 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_242
timestamp 1562078211
transform 1 0 23368 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_254
timestamp 1562078211
transform 1 0 24472 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_63_266
timestamp 1
transform 1 0 25576 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_274
timestamp 1
transform 1 0 26312 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_276
timestamp 1
transform 1 0 26496 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_297
timestamp 1
transform 1 0 28428 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_3
timestamp 1562078211
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_15
timestamp 1562078211
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_29
timestamp 1562078211
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_41
timestamp 1562078211
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_53
timestamp 1562078211
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_65
timestamp 1
transform 1 0 7084 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_91
timestamp 1
transform 1 0 9476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_95
timestamp 1
transform 1 0 9844 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_97
timestamp 1
transform 1 0 10028 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_136
timestamp 1
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_141
timestamp 1562078211
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_153
timestamp 1562078211
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_165
timestamp 1562078211
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_177
timestamp 1562078211
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_64_189
timestamp 1
transform 1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_193
timestamp 1
transform 1 0 18860 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_197
timestamp 1562078211
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_209
timestamp 1562078211
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_221
timestamp 1562078211
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_233
timestamp 1
transform 1 0 22540 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_235
timestamp 1
transform 1 0 22724 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_256
timestamp 1562078211
transform 1 0 24656 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_64_268
timestamp 1
transform 1 0 25760 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_276
timestamp 1
transform 1 0 26496 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_286
timestamp 1
transform 1 0 27416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_290
timestamp 1
transform 1 0 27784 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_3
timestamp 1562078211
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_15
timestamp 1562078211
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_27
timestamp 1562078211
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_39
timestamp 1562078211
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_65_51
timestamp 1
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_57
timestamp 1562078211
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_69
timestamp 1562078211
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_89
timestamp 1
transform 1 0 9292 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_65_98
timestamp 1
transform 1 0 10120 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_102
timestamp 1
transform 1 0 10488 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_65_113
timestamp 1
transform 1 0 11500 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_117
timestamp 1
transform 1 0 11868 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_119
timestamp 1
transform 1 0 12052 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_65_134
timestamp 1
transform 1 0 13432 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_138
timestamp 1
transform 1 0 13800 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_147
timestamp 1562078211
transform 1 0 14628 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_65_159
timestamp 1
transform 1 0 15732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_171
timestamp 1
transform 1 0 16836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_177
timestamp 1562078211
transform 1 0 17388 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_189
timestamp 1562078211
transform 1 0 18492 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_201
timestamp 1562078211
transform 1 0 19596 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_65_213
timestamp 1
transform 1 0 20700 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_221
timestamp 1
transform 1 0 21436 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_225
timestamp 1562078211
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_65_237
timestamp 1
transform 1 0 22908 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_250
timestamp 1562078211
transform 1 0 24104 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_262
timestamp 1562078211
transform 1 0 25208 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_65_274
timestamp 1
transform 1 0 26312 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_65_288
timestamp 1
transform 1 0 27600 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_296
timestamp 1
transform 1 0 28336 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_298
timestamp 1
transform 1 0 28520 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_3
timestamp 1562078211
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_15
timestamp 1562078211
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_29
timestamp 1562078211
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_41
timestamp 1562078211
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_53
timestamp 1562078211
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_66_65
timestamp 1
transform 1 0 7084 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_73
timestamp 1
transform 1 0 7820 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_75
timestamp 1
transform 1 0 8004 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_81
timestamp 1
transform 1 0 8556 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_66_85
timestamp 1
transform 1 0 8924 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_89
timestamp 1
transform 1 0 9292 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_112
timestamp 1562078211
transform 1 0 11408 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_66_124
timestamp 1
transform 1 0 12512 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_132
timestamp 1
transform 1 0 13248 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_141
timestamp 1
transform 1 0 14076 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_159
timestamp 1
transform 1 0 15732 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_167
timestamp 1
transform 1 0 16468 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_66_189
timestamp 1
transform 1 0 18492 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_193
timestamp 1
transform 1 0 18860 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_197
timestamp 1
transform 1 0 19228 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_208
timestamp 1
transform 1 0 20240 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_212
timestamp 1562078211
transform 1 0 20608 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_224
timestamp 1562078211
transform 1 0 21712 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_236
timestamp 1562078211
transform 1 0 22816 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_66_248
timestamp 1
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_253
timestamp 1562078211
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_265
timestamp 1562078211
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_277
timestamp 1
transform 1 0 26588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_285
timestamp 1562078211
transform 1 0 27324 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_297
timestamp 1
transform 1 0 28428 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_3
timestamp 1562078211
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_15
timestamp 1562078211
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_27
timestamp 1562078211
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_39
timestamp 1562078211
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_67_51
timestamp 1
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_57
timestamp 1562078211
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_69
timestamp 1
transform 1 0 7452 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_67_87
timestamp 1
transform 1 0 9108 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_91
timestamp 1
transform 1 0 9476 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_108
timestamp 1
transform 1 0 11040 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_113
timestamp 1562078211
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_67_125
timestamp 1
transform 1 0 12604 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_129
timestamp 1
transform 1 0 12972 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_67_136
timestamp 1
transform 1 0 13616 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_144
timestamp 1
transform 1 0 14352 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_149
timestamp 1562078211
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_161
timestamp 1
transform 1 0 15916 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_194
timestamp 1
transform 1 0 18952 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_220
timestamp 1
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_225
timestamp 1562078211
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_237
timestamp 1
transform 1 0 22908 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_245
timestamp 1562078211
transform 1 0 23644 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_257
timestamp 1562078211
transform 1 0 24748 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_67_269
timestamp 1
transform 1 0 25852 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_277
timestamp 1
transform 1 0 26588 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_281
timestamp 1562078211
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_67_293
timestamp 1
transform 1 0 28060 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_297
timestamp 1
transform 1 0 28428 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_3
timestamp 1562078211
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_15
timestamp 1562078211
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_29
timestamp 1562078211
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_41
timestamp 1562078211
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_53
timestamp 1562078211
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_65
timestamp 1562078211
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_77
timestamp 1
transform 1 0 8188 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_101
timestamp 1
transform 1 0 10396 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_122
timestamp 1
transform 1 0 12328 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_141
timestamp 1562078211
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_153
timestamp 1562078211
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_68_165
timestamp 1
transform 1 0 16284 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_189
timestamp 1
transform 1 0 18492 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_193
timestamp 1
transform 1 0 18860 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_226
timestamp 1562078211
transform 1 0 21896 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_68_238
timestamp 1
transform 1 0 23000 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_242
timestamp 1
transform 1 0 23368 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_258
timestamp 1562078211
transform 1 0 24840 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_270
timestamp 1562078211
transform 1 0 25944 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_282
timestamp 1562078211
transform 1 0 27048 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_68_294
timestamp 1
transform 1 0 28152 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_298
timestamp 1
transform 1 0 28520 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_3
timestamp 1562078211
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_15
timestamp 1562078211
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_27
timestamp 1562078211
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_39
timestamp 1562078211
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_69_51
timestamp 1
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_57
timestamp 1562078211
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_69
timestamp 1562078211
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_81
timestamp 1
transform 1 0 8556 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_69_91
timestamp 1
transform 1 0 9476 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_99
timestamp 1
transform 1 0 10212 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_101
timestamp 1
transform 1 0 10396 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_108
timestamp 1
transform 1 0 11040 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_113
timestamp 1
transform 1 0 11500 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_117
timestamp 1
transform 1 0 11868 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_135
timestamp 1562078211
transform 1 0 13524 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_147
timestamp 1562078211
transform 1 0 14628 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_69_159
timestamp 1
transform 1 0 15732 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_169
timestamp 1562078211
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_181
timestamp 1562078211
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_69_193
timestamp 1
transform 1 0 18860 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_201
timestamp 1
transform 1 0 19596 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_69_206
timestamp 1
transform 1 0 20056 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_220
timestamp 1
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_225
timestamp 1562078211
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_237
timestamp 1
transform 1 0 22908 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_239
timestamp 1
transform 1 0 23092 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_259
timestamp 1562078211
transform 1 0 24932 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_69_271
timestamp 1
transform 1 0 26036 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_292
timestamp 1
transform 1 0 27968 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_296
timestamp 1
transform 1 0 28336 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_298
timestamp 1
transform 1 0 28520 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_3
timestamp 1562078211
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_15
timestamp 1562078211
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_29
timestamp 1562078211
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_41
timestamp 1562078211
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_53
timestamp 1562078211
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_65
timestamp 1562078211
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_77
timestamp 1
transform 1 0 8188 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_81
timestamp 1
transform 1 0 8556 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_85
timestamp 1562078211
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_97
timestamp 1562078211
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_109
timestamp 1562078211
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_121
timestamp 1562078211
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_133
timestamp 1
transform 1 0 13340 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_137
timestamp 1
transform 1 0 13708 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_141
timestamp 1562078211
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_153
timestamp 1562078211
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_165
timestamp 1562078211
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_177
timestamp 1562078211
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_189
timestamp 1
transform 1 0 18492 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_193
timestamp 1
transform 1 0 18860 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_197
timestamp 1562078211
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_209
timestamp 1
transform 1 0 20332 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_219
timestamp 1562078211
transform 1 0 21252 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_231
timestamp 1
transform 1 0 22356 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_233
timestamp 1
transform 1 0 22540 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_70_248
timestamp 1
transform 1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_256
timestamp 1562078211
transform 1 0 24656 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_268
timestamp 1
transform 1 0 25760 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_70_293
timestamp 1
transform 1 0 28060 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_297
timestamp 1
transform 1 0 28428 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_3
timestamp 1562078211
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_15
timestamp 1562078211
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_27
timestamp 1562078211
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_39
timestamp 1562078211
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_51
timestamp 1
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_57
timestamp 1562078211
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_69
timestamp 1562078211
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_81
timestamp 1562078211
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_93
timestamp 1562078211
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_105
timestamp 1
transform 1 0 10764 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_109
timestamp 1
transform 1 0 11132 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_113
timestamp 1562078211
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_125
timestamp 1562078211
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_137
timestamp 1562078211
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_149
timestamp 1562078211
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_161
timestamp 1
transform 1 0 15916 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_165
timestamp 1
transform 1 0 16284 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_179
timestamp 1562078211
transform 1 0 17572 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_191
timestamp 1562078211
transform 1 0 18676 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_203
timestamp 1562078211
transform 1 0 19780 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_71_215
timestamp 1
transform 1 0 20884 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_225
timestamp 1562078211
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_237
timestamp 1
transform 1 0 22908 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_241
timestamp 1
transform 1 0 23276 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_245
timestamp 1
transform 1 0 23644 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_255
timestamp 1562078211
transform 1 0 24564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_267
timestamp 1
transform 1 0 25668 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_271
timestamp 1
transform 1 0 26036 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_297
timestamp 1
transform 1 0 28428 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_3
timestamp 1562078211
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_15
timestamp 1562078211
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_29
timestamp 1562078211
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_41
timestamp 1562078211
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_53
timestamp 1562078211
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_65
timestamp 1562078211
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_72_77
timestamp 1
transform 1 0 8188 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_81
timestamp 1
transform 1 0 8556 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_85
timestamp 1562078211
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_97
timestamp 1562078211
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_109
timestamp 1562078211
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_121
timestamp 1562078211
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_72_133
timestamp 1
transform 1 0 13340 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_137
timestamp 1
transform 1 0 13708 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_141
timestamp 1562078211
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_72_153
timestamp 1
transform 1 0 15180 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_157
timestamp 1
transform 1 0 15548 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_175
timestamp 1562078211
transform 1 0 17204 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_72_187
timestamp 1
transform 1 0 18308 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_197
timestamp 1
transform 1 0 19228 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_205
timestamp 1
transform 1 0 19964 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_215
timestamp 1562078211
transform 1 0 20884 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_72_227
timestamp 1
transform 1 0 21988 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_235
timestamp 1
transform 1 0 22724 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_253
timestamp 1562078211
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_265
timestamp 1562078211
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_280
timestamp 1562078211
transform 1 0 26864 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_72_292
timestamp 1
transform 1 0 27968 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_296
timestamp 1
transform 1 0 28336 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_298
timestamp 1
transform 1 0 28520 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_3
timestamp 1562078211
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_15
timestamp 1562078211
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_27
timestamp 1562078211
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_39
timestamp 1562078211
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_51
timestamp 1
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_57
timestamp 1562078211
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_69
timestamp 1562078211
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_81
timestamp 1562078211
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_93
timestamp 1562078211
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_105
timestamp 1
transform 1 0 10764 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_109
timestamp 1
transform 1 0 11132 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_113
timestamp 1
transform 1 0 11500 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_121
timestamp 1
transform 1 0 12236 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_123
timestamp 1
transform 1 0 12420 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_132
timestamp 1562078211
transform 1 0 13248 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_144
timestamp 1562078211
transform 1 0 14352 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_156
timestamp 1562078211
transform 1 0 15456 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_169
timestamp 1562078211
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_181
timestamp 1562078211
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_193
timestamp 1562078211
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_205
timestamp 1562078211
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_217
timestamp 1
transform 1 0 21068 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_221
timestamp 1
transform 1 0 21436 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_225
timestamp 1562078211
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_237
timestamp 1562078211
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_249
timestamp 1562078211
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_261
timestamp 1562078211
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_273
timestamp 1
transform 1 0 26220 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_277
timestamp 1
transform 1 0 26588 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_281
timestamp 1562078211
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_293
timestamp 1
transform 1 0 28060 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_297
timestamp 1
transform 1 0 28428 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_3
timestamp 1562078211
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_15
timestamp 1562078211
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_29
timestamp 1562078211
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_41
timestamp 1562078211
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_53
timestamp 1562078211
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_65
timestamp 1562078211
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_74_77
timestamp 1
transform 1 0 8188 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_81
timestamp 1
transform 1 0 8556 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_85
timestamp 1562078211
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_74_97
timestamp 1
transform 1 0 10028 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_105
timestamp 1
transform 1 0 10764 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_107
timestamp 1
transform 1 0 10948 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_74_135
timestamp 1
transform 1 0 13524 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_141
timestamp 1562078211
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_153
timestamp 1562078211
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_165
timestamp 1562078211
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_177
timestamp 1562078211
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_74_189
timestamp 1
transform 1 0 18492 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_193
timestamp 1
transform 1 0 18860 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_197
timestamp 1562078211
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_74_209
timestamp 1
transform 1 0 20332 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_225
timestamp 1562078211
transform 1 0 21804 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_237
timestamp 1562078211
transform 1 0 22908 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_249
timestamp 1
transform 1 0 24012 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_253
timestamp 1562078211
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_265
timestamp 1562078211
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_277
timestamp 1562078211
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_74_289
timestamp 1
transform 1 0 27692 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_297
timestamp 1
transform 1 0 28428 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_3
timestamp 1562078211
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_15
timestamp 1562078211
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_27
timestamp 1562078211
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_39
timestamp 1562078211
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_51
timestamp 1
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_57
timestamp 1562078211
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_69
timestamp 1562078211
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_81
timestamp 1562078211
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_93
timestamp 1562078211
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_105
timestamp 1
transform 1 0 10764 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_109
timestamp 1
transform 1 0 11132 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_142
timestamp 1562078211
transform 1 0 14168 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_154
timestamp 1562078211
transform 1 0 15272 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_166
timestamp 1
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_169
timestamp 1562078211
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_181
timestamp 1562078211
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_75_193
timestamp 1
transform 1 0 18860 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_201
timestamp 1
transform 1 0 19596 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_203
timestamp 1
transform 1 0 19780 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_75_220
timestamp 1
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_225
timestamp 1562078211
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_237
timestamp 1562078211
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_249
timestamp 1562078211
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_261
timestamp 1562078211
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_273
timestamp 1
transform 1 0 26220 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_277
timestamp 1
transform 1 0 26588 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_281
timestamp 1562078211
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_293
timestamp 1
transform 1 0 28060 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_297
timestamp 1
transform 1 0 28428 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_3
timestamp 1562078211
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_15
timestamp 1562078211
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_29
timestamp 1562078211
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_41
timestamp 1562078211
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_53
timestamp 1562078211
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_65
timestamp 1562078211
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_76_77
timestamp 1
transform 1 0 8188 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_81
timestamp 1
transform 1 0 8556 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_85
timestamp 1
transform 1 0 8924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_87
timestamp 1
transform 1 0 9108 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_104
timestamp 1
transform 1 0 10672 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_112
timestamp 1
transform 1 0 11408 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_149
timestamp 1562078211
transform 1 0 14812 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_161
timestamp 1562078211
transform 1 0 15916 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_173
timestamp 1562078211
transform 1 0 17020 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_76_185
timestamp 1
transform 1 0 18124 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_193
timestamp 1
transform 1 0 18860 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_197
timestamp 1562078211
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_209
timestamp 1562078211
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_221
timestamp 1562078211
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_233
timestamp 1562078211
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_76_245
timestamp 1
transform 1 0 23644 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_249
timestamp 1
transform 1 0 24012 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_253
timestamp 1562078211
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_265
timestamp 1562078211
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_277
timestamp 1562078211
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_76_289
timestamp 1
transform 1 0 27692 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_297
timestamp 1
transform 1 0 28428 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_3
timestamp 1562078211
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_15
timestamp 1562078211
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_27
timestamp 1562078211
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_39
timestamp 1562078211
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_77_51
timestamp 1
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_57
timestamp 1562078211
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_77_69
timestamp 1
transform 1 0 7452 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_113
timestamp 1
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_115
timestamp 1
transform 1 0 11684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_147
timestamp 1562078211
transform 1 0 14628 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_77_159
timestamp 1
transform 1 0 15732 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_169
timestamp 1562078211
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_181
timestamp 1562078211
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_193
timestamp 1562078211
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_205
timestamp 1562078211
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_77_217
timestamp 1
transform 1 0 21068 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_221
timestamp 1
transform 1 0 21436 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_225
timestamp 1562078211
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_237
timestamp 1562078211
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_249
timestamp 1562078211
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_261
timestamp 1562078211
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_77_273
timestamp 1
transform 1 0 26220 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_277
timestamp 1
transform 1 0 26588 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_281
timestamp 1562078211
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_77_293
timestamp 1
transform 1 0 28060 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_297
timestamp 1
transform 1 0 28428 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_3
timestamp 1562078211
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_15
timestamp 1562078211
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_29
timestamp 1562078211
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_41
timestamp 1562078211
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_53
timestamp 1562078211
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_65
timestamp 1
transform 1 0 7084 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_67
timestamp 1
transform 1 0 7268 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_78_93
timestamp 1
transform 1 0 9660 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_97
timestamp 1
transform 1 0 10028 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_123
timestamp 1
transform 1 0 12420 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_141
timestamp 1
transform 1 0 14076 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_155
timestamp 1562078211
transform 1 0 15364 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_167
timestamp 1562078211
transform 1 0 16468 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_179
timestamp 1562078211
transform 1 0 17572 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_78_191
timestamp 1
transform 1 0 18676 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_197
timestamp 1562078211
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_209
timestamp 1562078211
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_221
timestamp 1562078211
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_233
timestamp 1562078211
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_78_245
timestamp 1
transform 1 0 23644 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_249
timestamp 1
transform 1 0 24012 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_253
timestamp 1562078211
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_265
timestamp 1562078211
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_277
timestamp 1562078211
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_78_289
timestamp 1
transform 1 0 27692 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_297
timestamp 1
transform 1 0 28428 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_3
timestamp 1562078211
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_15
timestamp 1562078211
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_27
timestamp 1562078211
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_39
timestamp 1562078211
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_79_51
timestamp 1
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_79_57
timestamp 1
transform 1 0 6348 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_61
timestamp 1
transform 1 0 6716 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_68
timestamp 1562078211
transform 1 0 7360 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_80
timestamp 1562078211
transform 1 0 8464 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_92
timestamp 1562078211
transform 1 0 9568 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_79_104
timestamp 1
transform 1 0 10672 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_113
timestamp 1
transform 1 0 11500 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_117
timestamp 1
transform 1 0 11868 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_124
timestamp 1562078211
transform 1 0 12512 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_136
timestamp 1562078211
transform 1 0 13616 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_148
timestamp 1562078211
transform 1 0 14720 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_79_160
timestamp 1
transform 1 0 15824 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_169
timestamp 1562078211
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_181
timestamp 1562078211
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_193
timestamp 1562078211
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_205
timestamp 1562078211
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_79_217
timestamp 1
transform 1 0 21068 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_221
timestamp 1
transform 1 0 21436 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_225
timestamp 1562078211
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_237
timestamp 1562078211
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_249
timestamp 1562078211
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_261
timestamp 1562078211
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_79_273
timestamp 1
transform 1 0 26220 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_277
timestamp 1
transform 1 0 26588 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_281
timestamp 1562078211
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_79_293
timestamp 1
transform 1 0 28060 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_297
timestamp 1
transform 1 0 28428 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_3
timestamp 1562078211
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_15
timestamp 1562078211
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_29
timestamp 1562078211
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_41
timestamp 1562078211
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_53
timestamp 1562078211
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_65
timestamp 1562078211
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_77
timestamp 1
transform 1 0 8188 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_81
timestamp 1
transform 1 0 8556 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_85
timestamp 1562078211
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_97
timestamp 1562078211
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_109
timestamp 1562078211
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_121
timestamp 1562078211
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_133
timestamp 1
transform 1 0 13340 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_137
timestamp 1
transform 1 0 13708 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_141
timestamp 1562078211
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_153
timestamp 1562078211
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_165
timestamp 1562078211
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_177
timestamp 1562078211
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_189
timestamp 1
transform 1 0 18492 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_193
timestamp 1
transform 1 0 18860 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_197
timestamp 1562078211
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_209
timestamp 1562078211
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_221
timestamp 1562078211
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_233
timestamp 1562078211
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_245
timestamp 1
transform 1 0 23644 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_249
timestamp 1
transform 1 0 24012 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_253
timestamp 1562078211
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_265
timestamp 1562078211
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_277
timestamp 1562078211
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_80_289
timestamp 1
transform 1 0 27692 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_297
timestamp 1
transform 1 0 28428 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_3
timestamp 1562078211
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_15
timestamp 1562078211
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_27
timestamp 1562078211
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_39
timestamp 1562078211
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_51
timestamp 1
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_57
timestamp 1562078211
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_69
timestamp 1562078211
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_81
timestamp 1562078211
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_93
timestamp 1562078211
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_105
timestamp 1
transform 1 0 10764 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_109
timestamp 1
transform 1 0 11132 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_113
timestamp 1562078211
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_125
timestamp 1562078211
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_137
timestamp 1562078211
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_149
timestamp 1562078211
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_161
timestamp 1
transform 1 0 15916 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_165
timestamp 1
transform 1 0 16284 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_169
timestamp 1562078211
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_181
timestamp 1562078211
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_193
timestamp 1562078211
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_205
timestamp 1562078211
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_217
timestamp 1
transform 1 0 21068 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_221
timestamp 1
transform 1 0 21436 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_225
timestamp 1562078211
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_237
timestamp 1562078211
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_249
timestamp 1562078211
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_261
timestamp 1562078211
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_273
timestamp 1
transform 1 0 26220 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_277
timestamp 1
transform 1 0 26588 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_281
timestamp 1562078211
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_293
timestamp 1
transform 1 0 28060 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_297
timestamp 1
transform 1 0 28428 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_3
timestamp 1562078211
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_15
timestamp 1562078211
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_29
timestamp 1562078211
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_41
timestamp 1562078211
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_53
timestamp 1
transform 1 0 5980 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_55
timestamp 1
transform 1 0 6164 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_57
timestamp 1
transform 1 0 6348 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_62
timestamp 1562078211
transform 1 0 6808 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_82_74
timestamp 1
transform 1 0 7912 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_82
timestamp 1
transform 1 0 8648 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_85
timestamp 1562078211
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_97
timestamp 1562078211
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_109
timestamp 1
transform 1 0 11132 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_113
timestamp 1562078211
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_125
timestamp 1562078211
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_137
timestamp 1
transform 1 0 13708 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_141
timestamp 1562078211
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_153
timestamp 1562078211
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_165
timestamp 1
transform 1 0 16284 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_169
timestamp 1562078211
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_181
timestamp 1562078211
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_193
timestamp 1
transform 1 0 18860 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_197
timestamp 1562078211
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_209
timestamp 1562078211
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_221
timestamp 1
transform 1 0 21436 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_223
timestamp 1
transform 1 0 21620 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_225
timestamp 1562078211
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_237
timestamp 1562078211
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_249
timestamp 1
transform 1 0 24012 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_253
timestamp 1562078211
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_265
timestamp 1562078211
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_277
timestamp 1
transform 1 0 26588 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_279
timestamp 1
transform 1 0 26772 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_281
timestamp 1562078211
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_82_293
timestamp 1
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_297
timestamp 1
transform 1 0 28428 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform 1 0 11960 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 13248 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform 1 0 10396 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform 1 0 11040 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform 1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform 1 0 10120 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform 1 0 10396 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform 1 0 11132 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 10672 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 11316 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 12420 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform 1 0 11040 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform 1 0 6900 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 7176 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 12512 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 10120 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform 1 0 6900 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 11408 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 9476 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform 1 0 6532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 9292 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform 1 0 8648 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 8832 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 10396 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 6440 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 8556 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 6256 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform -1 0 9476 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform 1 0 14168 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 9568 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform -1 0 8188 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform -1 0 7084 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform -1 0 7636 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform -1 0 9660 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform -1 0 6532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform -1 0 14812 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform -1 0 9844 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 5612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform -1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform -1 0 6440 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform -1 0 9660 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform -1 0 7084 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform -1 0 19136 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform -1 0 18308 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform -1 0 16468 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform -1 0 21988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform -1 0 27416 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform 1 0 26128 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1
transform -1 0 28152 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1
transform -1 0 25116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1
transform -1 0 24012 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1
transform -1 0 20700 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1
transform 1 0 20884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1
transform -1 0 26496 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1
transform -1 0 25668 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1
transform -1 0 26680 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1
transform -1 0 28336 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1
transform -1 0 17388 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1
transform -1 0 20516 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1
transform -1 0 19780 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1
transform -1 0 28612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1
transform -1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1
transform -1 0 22908 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1
transform -1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1
transform 1 0 17020 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1
transform -1 0 26956 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1
transform -1 0 23828 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1
transform -1 0 21068 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1
transform -1 0 21252 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1
transform 1 0 20792 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1
transform -1 0 14720 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1
transform -1 0 17480 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1
transform -1 0 20332 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1
transform 1 0 19228 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1
transform -1 0 21804 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform -1 0 1656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 6808 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1656 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform 1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap19
timestamp 1
transform -1 0 12420 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1
transform 1 0 28244 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1
transform 1 0 28244 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform 1 0 28244 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_83
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_84
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_85
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_86
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_87
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_88
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_89
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_90
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_91
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_92
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_93
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_94
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_95
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_96
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_97
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_98
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_99
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_100
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_101
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_102
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_103
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_104
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_105
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_106
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_107
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_108
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_109
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_110
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_111
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_112
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_113
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_114
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_115
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_116
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_117
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_118
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_119
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_120
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_121
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_122
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_123
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_124
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_125
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_126
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_127
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_128
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_129
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_130
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_131
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_132
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_133
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_134
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_135
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_136
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_137
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1
transform -1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_138
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1
transform -1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_139
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1
transform -1 0 28888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_140
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1
transform -1 0 28888 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_141
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1
transform -1 0 28888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_142
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1
transform -1 0 28888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_143
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1
transform -1 0 28888 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_144
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1
transform -1 0 28888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_145
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1
transform -1 0 28888 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_146
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1
transform -1 0 28888 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_147
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1
transform -1 0 28888 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_148
timestamp 1
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1
transform -1 0 28888 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_149
timestamp 1
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1
transform -1 0 28888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_150
timestamp 1
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1
transform -1 0 28888 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_151
timestamp 1
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1
transform -1 0 28888 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_152
timestamp 1
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 1
transform -1 0 28888 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_153
timestamp 1
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 1
transform -1 0 28888 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_154
timestamp 1
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 1
transform -1 0 28888 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_155
timestamp 1
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 1
transform -1 0 28888 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_156
timestamp 1
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 1
transform -1 0 28888 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_157
timestamp 1
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 1
transform -1 0 28888 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_158
timestamp 1
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 1
transform -1 0 28888 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_159
timestamp 1
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 1
transform -1 0 28888 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_160
timestamp 1
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 1
transform -1 0 28888 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_161
timestamp 1
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 1
transform -1 0 28888 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_162
timestamp 1
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 1
transform -1 0 28888 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_163
timestamp 1
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 1
transform -1 0 28888 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_164
timestamp 1
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 1
transform -1 0 28888 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_165
timestamp 1
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 1
transform -1 0 28888 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_34
timestamp 1
transform 1 0 28336 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_35
timestamp 1
transform -1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_36
timestamp 1
transform 1 0 28336 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_37
timestamp 1
transform -1 0 1656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_38
timestamp 1
transform -1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_39
timestamp 1
transform -1 0 1656 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_40
timestamp 1
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_41
timestamp 1
transform 1 0 27968 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_42
timestamp 1
transform -1 0 1656 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_43
timestamp 1
transform -1 0 28612 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_166
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_167
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_168
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_169
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_170
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_171
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_172
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_173
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_174
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_175
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_176
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_177
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_178
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_179
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_180
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_181
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_182
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_183
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_184
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_185
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_186
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_187
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_188
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_189
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_190
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_191
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_192
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_193
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_194
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_195
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_196
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_197
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_198
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_199
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_200
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_201
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_202
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_203
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_204
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_205
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_206
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_207
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_208
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_209
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_210
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_211
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_212
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_213
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_214
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_215
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_216
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_217
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_218
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_219
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_220
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_221
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_222
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_223
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_224
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_225
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_226
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_227
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_228
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_229
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_230
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_231
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_232
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_233
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_234
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_235
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_236
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_237
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_238
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_239
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_240
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_241
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_242
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_243
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_244
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_245
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_246
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_247
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_248
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_249
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_250
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_251
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_252
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_253
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_254
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_255
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_256
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_257
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_258
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_259
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_260
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_261
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_262
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_263
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_264
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_265
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_266
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_267
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_268
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_269
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_270
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_271
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_272
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_273
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_274
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_275
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_276
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_277
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_278
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_279
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_280
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_281
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_282
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_283
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_284
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_285
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_286
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_287
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_288
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_289
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_290
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_291
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_292
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_293
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_294
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_295
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_296
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_297
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_298
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_299
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_300
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_301
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_302
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_303
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_304
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_305
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_306
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_307
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_308
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_309
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_310
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_311
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_312
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_313
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_314
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_315
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_316
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_317
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_318
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_319
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_320
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_321
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_322
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_323
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_324
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_325
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_326
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_327
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_328
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_329
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_330
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_331
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_332
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_333
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_334
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_335
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_336
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_337
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_338
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_339
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_340
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_341
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_342
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_343
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_344
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_345
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_346
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_347
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_348
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_349
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_350
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_351
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_352
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_353
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_354
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_355
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_356
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_357
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_358
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_359
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_360
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_361
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_362
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_363
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_364
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_365
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_366
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_367
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_368
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_369
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_370
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_371
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_372
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_373
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_374
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_375
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_376
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_377
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_378
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_379
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_380
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_381
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_382
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_383
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_384
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_385
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_386
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_387
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_388
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_389
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_390
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_391
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_392
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_393
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_394
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_395
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_396
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_397
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_398
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_399
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_400
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_401
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_402
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_403
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_404
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_405
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_406
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_407
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_408
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_409
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_410
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_411
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_412
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_413
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_414
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_415
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_416
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_417
timestamp 1
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_418
timestamp 1
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_419
timestamp 1
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_420
timestamp 1
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_421
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_422
timestamp 1
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_423
timestamp 1
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_424
timestamp 1
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_425
timestamp 1
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_426
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_427
timestamp 1
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_428
timestamp 1
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_429
timestamp 1
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_430
timestamp 1
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_431
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_432
timestamp 1
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_433
timestamp 1
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_434
timestamp 1
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_435
timestamp 1
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_436
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_437
timestamp 1
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_438
timestamp 1
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_439
timestamp 1
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_440
timestamp 1
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_441
timestamp 1
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_442
timestamp 1
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_443
timestamp 1
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_444
timestamp 1
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_445
timestamp 1
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_446
timestamp 1
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_447
timestamp 1
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_448
timestamp 1
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_449
timestamp 1
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_450
timestamp 1
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_451
timestamp 1
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_452
timestamp 1
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_453
timestamp 1
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_454
timestamp 1
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_455
timestamp 1
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_456
timestamp 1
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_457
timestamp 1
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_458
timestamp 1
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_459
timestamp 1
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_460
timestamp 1
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_461
timestamp 1
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_462
timestamp 1
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_463
timestamp 1
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_464
timestamp 1
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_465
timestamp 1
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_466
timestamp 1
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_467
timestamp 1
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_468
timestamp 1
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_469
timestamp 1
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_470
timestamp 1
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_471
timestamp 1
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_472
timestamp 1
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_473
timestamp 1
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_474
timestamp 1
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_475
timestamp 1
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_476
timestamp 1
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_477
timestamp 1
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_478
timestamp 1
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_479
timestamp 1
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_480
timestamp 1
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_481
timestamp 1
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_482
timestamp 1
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_483
timestamp 1
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_484
timestamp 1
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_485
timestamp 1
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_486
timestamp 1
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_487
timestamp 1
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_488
timestamp 1
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_489
timestamp 1
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_490
timestamp 1
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_491
timestamp 1
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_492
timestamp 1
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_493
timestamp 1
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_494
timestamp 1
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_495
timestamp 1
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_496
timestamp 1
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_497
timestamp 1
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_498
timestamp 1
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_499
timestamp 1
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_500
timestamp 1
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_501
timestamp 1
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_502
timestamp 1
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_503
timestamp 1
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_504
timestamp 1
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_505
timestamp 1
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_506
timestamp 1
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_507
timestamp 1
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_508
timestamp 1
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_509
timestamp 1
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_510
timestamp 1
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_511
timestamp 1
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_512
timestamp 1
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_513
timestamp 1
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_514
timestamp 1
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_515
timestamp 1
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_516
timestamp 1
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_517
timestamp 1
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_518
timestamp 1
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_519
timestamp 1
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_520
timestamp 1
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_521
timestamp 1
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_522
timestamp 1
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_523
timestamp 1
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_524
timestamp 1
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_525
timestamp 1
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_526
timestamp 1
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_527
timestamp 1
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_528
timestamp 1
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_529
timestamp 1
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_530
timestamp 1
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_531
timestamp 1
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_532
timestamp 1
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_533
timestamp 1
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_534
timestamp 1
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_535
timestamp 1
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_536
timestamp 1
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_537
timestamp 1
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_538
timestamp 1
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_539
timestamp 1
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_540
timestamp 1
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_541
timestamp 1
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_542
timestamp 1
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_543
timestamp 1
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_544
timestamp 1
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_545
timestamp 1
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_546
timestamp 1
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_547
timestamp 1
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_548
timestamp 1
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_549
timestamp 1
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_550
timestamp 1
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_551
timestamp 1
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_552
timestamp 1
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_553
timestamp 1
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_554
timestamp 1
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_555
timestamp 1
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_556
timestamp 1
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_557
timestamp 1
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_558
timestamp 1
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_559
timestamp 1
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_560
timestamp 1
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_561
timestamp 1
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_562
timestamp 1
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_563
timestamp 1
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_564
timestamp 1
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_565
timestamp 1
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_566
timestamp 1
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_567
timestamp 1
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_568
timestamp 1
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_569
timestamp 1
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_570
timestamp 1
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_571
timestamp 1
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_572
timestamp 1
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_573
timestamp 1
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_574
timestamp 1
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_575
timestamp 1
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_576
timestamp 1
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_577
timestamp 1
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_578
timestamp 1
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_579
timestamp 1
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_580
timestamp 1
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_581
timestamp 1
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_582
timestamp 1
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_583
timestamp 1
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_584
timestamp 1
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_585
timestamp 1
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_586
timestamp 1
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_587
timestamp 1
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_588
timestamp 1
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_589
timestamp 1
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_590
timestamp 1
transform 1 0 26864 0 1 46784
box -38 -48 130 592
<< labels >>
flabel metal2 s 24490 49200 24546 50000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 enc0_a
port 1 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 enc0_b
port 2 nsew signal input
flabel metal2 s 6458 49200 6514 50000 0 FreeSans 224 90 0 0 enc1_a
port 3 nsew signal input
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 enc1_b
port 4 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 enc2_a
port 5 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 enc2_b
port 6 nsew signal input
flabel metal3 s 29200 22448 30000 22568 0 FreeSans 480 0 0 0 io_oeb_high[0]
port 7 nsew signal output
flabel metal3 s 29200 19728 30000 19848 0 FreeSans 480 0 0 0 io_oeb_high[1]
port 8 nsew signal output
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 io_oeb_high[2]
port 9 nsew signal output
flabel metal3 s 29200 27888 30000 28008 0 FreeSans 480 0 0 0 io_oeb_high[3]
port 10 nsew signal output
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 io_oeb_high[4]
port 11 nsew signal output
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 io_oeb_high[5]
port 12 nsew signal output
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 io_oeb_low[0]
port 13 nsew signal output
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 io_oeb_low[1]
port 14 nsew signal output
flabel metal3 s 29200 15648 30000 15768 0 FreeSans 480 0 0 0 io_oeb_low[2]
port 15 nsew signal output
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 io_oeb_low[3]
port 16 nsew signal output
flabel metal3 s 29200 31288 30000 31408 0 FreeSans 480 0 0 0 pwm0_out
port 17 nsew signal output
flabel metal3 s 29200 35368 30000 35488 0 FreeSans 480 0 0 0 pwm1_out
port 18 nsew signal output
flabel metal3 s 29200 16328 30000 16448 0 FreeSans 480 0 0 0 pwm2_out
port 19 nsew signal output
flabel metal3 s 29200 8168 30000 8288 0 FreeSans 480 0 0 0 reset
port 20 nsew signal input
flabel metal3 s 29200 23128 30000 23248 0 FreeSans 480 0 0 0 sync
port 21 nsew signal output
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 22 nsew power bidirectional
flabel metal4 s 4868 2128 5188 47376 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
rlabel metal1 14996 47328 14996 47328 0 vccd1
rlabel metal1 14996 46784 14996 46784 0 vssd1
rlabel metal1 9092 27030 9092 27030 0 _000_
rlabel metal1 3710 29546 3710 29546 0 _001_
rlabel metal1 5285 30226 5285 30226 0 _002_
rlabel metal1 6021 29546 6021 29546 0 _003_
rlabel via1 6665 30294 6665 30294 0 _004_
rlabel metal1 8362 29546 8362 29546 0 _005_
rlabel metal1 8954 29206 8954 29206 0 _006_
rlabel metal1 10084 30226 10084 30226 0 _007_
rlabel metal2 8694 31586 8694 31586 0 _008_
rlabel metal2 7498 22780 7498 22780 0 _009_
rlabel viali 3445 24786 3445 24786 0 _010_
rlabel metal2 4830 24582 4830 24582 0 _011_
rlabel metal1 6693 23766 6693 23766 0 _012_
rlabel metal2 7866 24786 7866 24786 0 _013_
rlabel metal1 5653 23018 5653 23018 0 _014_
rlabel via1 5653 18734 5653 18734 0 _015_
rlabel metal1 5515 19346 5515 19346 0 _016_
rlabel metal2 6394 19618 6394 19618 0 _017_
rlabel metal1 13064 42194 13064 42194 0 _018_
rlabel metal1 7482 44778 7482 44778 0 _019_
rlabel metal1 9052 43758 9052 43758 0 _020_
rlabel metal1 9598 44438 9598 44438 0 _021_
rlabel metal2 11546 44370 11546 44370 0 _022_
rlabel via1 11357 42670 11357 42670 0 _023_
rlabel metal1 13064 42874 13064 42874 0 _024_
rlabel metal2 12650 44268 12650 44268 0 _025_
rlabel metal1 14408 44370 14408 44370 0 _026_
rlabel metal1 10948 36890 10948 36890 0 _027_
rlabel metal1 4186 33626 4186 33626 0 _028_
rlabel metal1 6946 35632 6946 35632 0 _029_
rlabel metal1 9476 35734 9476 35734 0 _030_
rlabel metal2 11914 35462 11914 35462 0 _031_
rlabel metal2 8050 37026 8050 37026 0 _032_
rlabel metal1 8050 38522 8050 38522 0 _033_
rlabel metal1 9000 39338 9000 39338 0 _034_
rlabel metal2 9890 38726 9890 38726 0 _035_
rlabel metal1 12282 10540 12282 10540 0 _036_
rlabel metal2 5658 8738 5658 8738 0 _037_
rlabel metal2 7314 9078 7314 9078 0 _038_
rlabel metal1 9338 10778 9338 10778 0 _039_
rlabel metal1 9517 11798 9517 11798 0 _040_
rlabel metal2 10994 10200 10994 10200 0 _041_
rlabel metal1 10457 7786 10457 7786 0 _042_
rlabel metal1 9747 8534 9747 8534 0 _043_
rlabel metal2 12190 9350 12190 9350 0 _044_
rlabel metal1 11500 16422 11500 16422 0 _045_
rlabel via1 16877 16558 16877 16558 0 _046_
rlabel metal1 17480 15470 17480 15470 0 _047_
rlabel metal1 18717 17238 18717 17238 0 _048_
rlabel metal2 19642 18258 19642 18258 0 _049_
rlabel metal1 20516 17306 20516 17306 0 _050_
rlabel metal1 22356 17850 22356 17850 0 _051_
rlabel metal1 23736 17306 23736 17306 0 _052_
rlabel metal1 25208 17850 25208 17850 0 _053_
rlabel metal1 9384 26010 9384 26010 0 _054_
rlabel metal2 3450 15844 3450 15844 0 _055_
rlabel metal1 6562 16150 6562 16150 0 _056_
rlabel metal1 6838 15402 6838 15402 0 _057_
rlabel metal1 7636 14586 7636 14586 0 _058_
rlabel metal2 9706 14790 9706 14790 0 _059_
rlabel metal1 11408 16762 11408 16762 0 _060_
rlabel metal1 9936 17510 9936 17510 0 _061_
rlabel metal2 9062 18530 9062 18530 0 _062_
rlabel metal1 14536 20026 14536 20026 0 _063_
rlabel metal1 12640 19822 12640 19822 0 _064_
rlabel via1 12277 26282 12277 26282 0 _065_
rlabel metal1 14572 26350 14572 26350 0 _066_
rlabel via1 11541 30702 11541 30702 0 _067_
rlabel metal2 13294 33286 13294 33286 0 _068_
rlabel metal2 16238 34374 16238 34374 0 _069_
rlabel metal1 16518 29614 16518 29614 0 _070_
rlabel metal1 13013 39338 13013 39338 0 _071_
rlabel metal1 6808 23086 6808 23086 0 _072_
rlabel metal2 16698 41378 16698 41378 0 _073_
rlabel metal1 16790 38896 16790 38896 0 _074_
rlabel metal2 19550 38760 19550 38760 0 _075_
rlabel metal2 20194 42534 20194 42534 0 _076_
rlabel metal2 23230 37026 23230 37026 0 _077_
rlabel metal1 23317 41514 23317 41514 0 _078_
rlabel metal1 26986 41174 26986 41174 0 _079_
rlabel metal1 26940 36822 26940 36822 0 _080_
rlabel metal2 12650 12818 12650 12818 0 _081_
rlabel metal1 12374 36890 12374 36890 0 _082_
rlabel metal2 14766 8738 14766 8738 0 _083_
rlabel metal2 15226 10438 15226 10438 0 _084_
rlabel via1 17245 8466 17245 8466 0 _085_
rlabel metal1 19448 7854 19448 7854 0 _086_
rlabel via1 22121 8534 22121 8534 0 _087_
rlabel metal2 22034 13022 22034 13022 0 _088_
rlabel metal1 24324 8942 24324 8942 0 _089_
rlabel metal1 24968 13294 24968 13294 0 _090_
rlabel metal2 27094 29614 27094 29614 0 _091_
rlabel metal1 10534 16626 10534 16626 0 _092_
rlabel metal2 26818 35122 26818 35122 0 _093_
rlabel metal1 15083 17578 15083 17578 0 _094_
rlabel metal2 15686 19618 15686 19618 0 _095_
rlabel via1 17162 21998 17162 21998 0 _096_
rlabel metal1 20198 22610 20198 22610 0 _097_
rlabel via1 18533 22610 18533 22610 0 _098_
rlabel metal1 19120 27370 19120 27370 0 _099_
rlabel metal2 22034 27812 22034 27812 0 _100_
rlabel metal2 21574 27200 21574 27200 0 _101_
rlabel metal1 26174 16660 26174 16660 0 _102_
rlabel metal1 17970 33558 17970 33558 0 _103_
rlabel metal2 19274 32572 19274 32572 0 _104_
rlabel via1 20750 32810 20750 32810 0 _105_
rlabel metal2 22126 33286 22126 33286 0 _106_
rlabel metal2 22218 32674 22218 32674 0 _107_
rlabel metal2 24426 32198 24426 32198 0 _108_
rlabel via1 25433 32402 25433 32402 0 _109_
rlabel metal1 27048 31994 27048 31994 0 _110_
rlabel metal1 24794 16082 24794 16082 0 _111_
rlabel metal1 24242 15946 24242 15946 0 _112_
rlabel metal2 22218 15538 22218 15538 0 _113_
rlabel metal1 19090 14382 19090 14382 0 _114_
rlabel metal1 18538 14382 18538 14382 0 _115_
rlabel metal2 17250 14722 17250 14722 0 _116_
rlabel metal2 16974 13566 16974 13566 0 _117_
rlabel metal1 27048 36890 27048 36890 0 _118_
rlabel metal2 27278 34204 27278 34204 0 _119_
rlabel via1 24334 34646 24334 34646 0 _120_
rlabel viali 23598 34578 23598 34578 0 _121_
rlabel metal1 21574 39338 21574 39338 0 _122_
rlabel metal1 20378 38182 20378 38182 0 _123_
rlabel metal1 17986 38250 17986 38250 0 _124_
rlabel metal2 18584 38930 18584 38930 0 _125_
rlabel metal1 17342 33626 17342 33626 0 _126_
rlabel metal1 13570 31790 13570 31790 0 _127_
rlabel metal2 17526 28016 17526 28016 0 _128_
rlabel metal1 15042 23630 15042 23630 0 _129_
rlabel metal2 15318 23222 15318 23222 0 _130_
rlabel metal1 12926 10710 12926 10710 0 _131_
rlabel metal1 9660 29138 9660 29138 0 _132_
rlabel metal2 8970 30124 8970 30124 0 _133_
rlabel metal1 9292 28526 9292 28526 0 _134_
rlabel metal1 10074 28458 10074 28458 0 _135_
rlabel metal1 7682 21998 7682 21998 0 _136_
rlabel metal2 6394 23188 6394 23188 0 _137_
rlabel metal2 7130 23290 7130 23290 0 _138_
rlabel metal2 7130 22542 7130 22542 0 _139_
rlabel metal1 12788 43962 12788 43962 0 _140_
rlabel metal2 12834 43146 12834 43146 0 _141_
rlabel metal1 12650 43826 12650 43826 0 _142_
rlabel metal1 12604 42670 12604 42670 0 _143_
rlabel metal1 9706 36754 9706 36754 0 _144_
rlabel metal1 10718 36720 10718 36720 0 _145_
rlabel metal1 10166 37128 10166 37128 0 _146_
rlabel metal1 10902 37094 10902 37094 0 _147_
rlabel metal1 10626 9690 10626 9690 0 _148_
rlabel metal1 11638 10234 11638 10234 0 _149_
rlabel metal1 10810 9146 10810 9146 0 _150_
rlabel metal2 10166 10472 10166 10472 0 _151_
rlabel metal2 10534 15198 10534 15198 0 _152_
rlabel metal1 10304 16218 10304 16218 0 _153_
rlabel metal1 11270 16694 11270 16694 0 _154_
rlabel metal2 10994 15300 10994 15300 0 _155_
rlabel metal1 17986 15504 17986 15504 0 _156_
rlabel metal1 18584 17646 18584 17646 0 _157_
rlabel metal1 21260 17306 21260 17306 0 _158_
rlabel metal2 20930 17952 20930 17952 0 _159_
rlabel metal1 19826 17680 19826 17680 0 _160_
rlabel metal1 23046 18768 23046 18768 0 _161_
rlabel metal2 20746 17918 20746 17918 0 _162_
rlabel metal2 23138 17884 23138 17884 0 _163_
rlabel metal1 22816 17306 22816 17306 0 _164_
rlabel metal1 23920 17850 23920 17850 0 _165_
rlabel metal2 23506 17884 23506 17884 0 _166_
rlabel metal2 25438 17340 25438 17340 0 _167_
rlabel metal2 11454 23324 11454 23324 0 _168_
rlabel metal2 11270 23290 11270 23290 0 _169_
rlabel metal2 10626 22916 10626 22916 0 _170_
rlabel metal1 12972 31858 12972 31858 0 _171_
rlabel metal2 14398 20026 14398 20026 0 _172_
rlabel metal1 11914 22984 11914 22984 0 _173_
rlabel metal2 11730 22780 11730 22780 0 _174_
rlabel metal1 13478 24786 13478 24786 0 _175_
rlabel metal2 12466 21794 12466 21794 0 _176_
rlabel metal1 13110 21862 13110 21862 0 _177_
rlabel metal2 12190 20842 12190 20842 0 _178_
rlabel metal2 12466 20604 12466 20604 0 _179_
rlabel metal2 13018 20604 13018 20604 0 _180_
rlabel metal2 12282 23596 12282 23596 0 _181_
rlabel metal1 12213 25874 12213 25874 0 _182_
rlabel metal2 12190 25500 12190 25500 0 _183_
rlabel metal1 13110 25466 13110 25466 0 _184_
rlabel metal1 12742 25908 12742 25908 0 _185_
rlabel metal2 13018 25636 13018 25636 0 _186_
rlabel metal2 13110 26282 13110 26282 0 _187_
rlabel metal2 13478 26724 13478 26724 0 _188_
rlabel metal2 14030 27132 14030 27132 0 _189_
rlabel metal1 14398 31858 14398 31858 0 _190_
rlabel metal1 14122 31790 14122 31790 0 _191_
rlabel metal1 13616 31994 13616 31994 0 _192_
rlabel metal1 13570 26554 13570 26554 0 _193_
rlabel metal2 12926 28900 12926 28900 0 _194_
rlabel metal1 12420 32334 12420 32334 0 _195_
rlabel metal1 12512 32402 12512 32402 0 _196_
rlabel metal2 12006 31756 12006 31756 0 _197_
rlabel metal1 13294 32300 13294 32300 0 _198_
rlabel metal1 12742 32844 12742 32844 0 _199_
rlabel metal1 14076 32266 14076 32266 0 _200_
rlabel metal1 12604 32946 12604 32946 0 _201_
rlabel metal1 15548 33558 15548 33558 0 _202_
rlabel metal1 15778 33354 15778 33354 0 _203_
rlabel metal1 15594 33456 15594 33456 0 _204_
rlabel metal1 13294 32402 13294 32402 0 _205_
rlabel metal2 15318 32708 15318 32708 0 _206_
rlabel metal1 15962 33592 15962 33592 0 _207_
rlabel metal2 16698 33796 16698 33796 0 _208_
rlabel metal1 15686 32742 15686 32742 0 _209_
rlabel metal2 15686 30464 15686 30464 0 _210_
rlabel metal1 15870 30294 15870 30294 0 _211_
rlabel metal1 16192 30090 16192 30090 0 _212_
rlabel metal1 15686 38352 15686 38352 0 _213_
rlabel metal1 15410 38182 15410 38182 0 _214_
rlabel metal2 15410 38522 15410 38522 0 _215_
rlabel metal1 17756 39338 17756 39338 0 _216_
rlabel metal1 16882 41038 16882 41038 0 _217_
rlabel metal1 17158 37672 17158 37672 0 _218_
rlabel metal1 17426 37978 17426 37978 0 _219_
rlabel metal1 17894 39372 17894 39372 0 _220_
rlabel metal1 16652 38318 16652 38318 0 _221_
rlabel metal1 18538 38250 18538 38250 0 _222_
rlabel metal1 17158 38318 17158 38318 0 _223_
rlabel metal2 16790 38998 16790 38998 0 _224_
rlabel metal1 17296 38386 17296 38386 0 _225_
rlabel metal2 16882 38794 16882 38794 0 _226_
rlabel metal2 19918 39168 19918 39168 0 _227_
rlabel metal2 20102 38964 20102 38964 0 _228_
rlabel metal1 20654 39610 20654 39610 0 _229_
rlabel metal2 19826 39610 19826 39610 0 _230_
rlabel metal1 20240 39066 20240 39066 0 _231_
rlabel metal1 19596 38318 19596 38318 0 _232_
rlabel metal2 21022 40324 21022 40324 0 _233_
rlabel metal1 21206 40528 21206 40528 0 _234_
rlabel metal2 21114 41072 21114 41072 0 _235_
rlabel metal1 20516 40698 20516 40698 0 _236_
rlabel metal1 20470 41718 20470 41718 0 _237_
rlabel metal1 23920 39610 23920 39610 0 _238_
rlabel metal1 24610 39372 24610 39372 0 _239_
rlabel metal2 23322 39474 23322 39474 0 _240_
rlabel metal2 20470 39644 20470 39644 0 _241_
rlabel metal2 23138 39066 23138 39066 0 _242_
rlabel metal1 23690 37978 23690 37978 0 _243_
rlabel metal2 23322 37196 23322 37196 0 _244_
rlabel metal1 23644 40358 23644 40358 0 _245_
rlabel metal1 23460 40154 23460 40154 0 _246_
rlabel metal2 23230 40868 23230 40868 0 _247_
rlabel metal1 23690 41106 23690 41106 0 _248_
rlabel metal1 27186 40494 27186 40494 0 _249_
rlabel metal2 27922 40256 27922 40256 0 _250_
rlabel metal1 26726 40154 26726 40154 0 _251_
rlabel metal1 24564 39950 24564 39950 0 _252_
rlabel metal1 26266 41038 26266 41038 0 _253_
rlabel metal2 27186 40732 27186 40732 0 _254_
rlabel metal1 26772 40698 26772 40698 0 _255_
rlabel metal1 27324 38318 27324 38318 0 _256_
rlabel metal1 27094 37978 27094 37978 0 _257_
rlabel metal2 27094 37706 27094 37706 0 _258_
rlabel metal1 27002 37366 27002 37366 0 _259_
rlabel metal1 14122 14858 14122 14858 0 _260_
rlabel metal1 14444 15062 14444 15062 0 _261_
rlabel metal1 14674 14960 14674 14960 0 _262_
rlabel metal1 15318 14790 15318 14790 0 _263_
rlabel metal2 14950 8908 14950 8908 0 _264_
rlabel metal2 15502 13804 15502 13804 0 _265_
rlabel metal2 15318 13770 15318 13770 0 _266_
rlabel metal1 16100 13362 16100 13362 0 _267_
rlabel metal1 15916 11322 15916 11322 0 _268_
rlabel metal1 16376 12886 16376 12886 0 _269_
rlabel metal1 16606 12818 16606 12818 0 _270_
rlabel metal2 15134 11356 15134 11356 0 _271_
rlabel metal1 15962 11220 15962 11220 0 _272_
rlabel metal1 15364 10030 15364 10030 0 _273_
rlabel metal1 17526 12682 17526 12682 0 _274_
rlabel metal2 18630 9758 18630 9758 0 _275_
rlabel metal2 18078 11084 18078 11084 0 _276_
rlabel metal2 18446 10268 18446 10268 0 _277_
rlabel metal1 17710 8942 17710 8942 0 _278_
rlabel metal1 19090 9622 19090 9622 0 _279_
rlabel metal1 19504 10506 19504 10506 0 _280_
rlabel metal2 19734 9452 19734 9452 0 _281_
rlabel metal2 18906 8636 18906 8636 0 _282_
rlabel metal1 21850 9554 21850 9554 0 _283_
rlabel metal2 19458 10132 19458 10132 0 _284_
rlabel metal1 21850 11152 21850 11152 0 _285_
rlabel metal2 22494 9146 22494 9146 0 _286_
rlabel metal2 21942 9010 21942 9010 0 _287_
rlabel metal1 21620 12206 21620 12206 0 _288_
rlabel metal1 21528 11322 21528 11322 0 _289_
rlabel metal1 21942 12104 21942 12104 0 _290_
rlabel metal1 21896 12410 21896 12410 0 _291_
rlabel metal2 24794 10438 24794 10438 0 _292_
rlabel metal1 25024 10710 25024 10710 0 _293_
rlabel metal1 24840 10030 24840 10030 0 _294_
rlabel metal2 22310 11662 22310 11662 0 _295_
rlabel metal2 24518 10914 24518 10914 0 _296_
rlabel metal1 25024 9690 25024 9690 0 _297_
rlabel metal1 23966 9520 23966 9520 0 _298_
rlabel metal1 25300 10778 25300 10778 0 _299_
rlabel metal1 25162 12716 25162 12716 0 _300_
rlabel metal1 25300 12954 25300 12954 0 _301_
rlabel metal1 24794 13498 24794 13498 0 _302_
rlabel metal2 18446 28934 18446 28934 0 _303_
rlabel metal2 17710 27234 17710 27234 0 _304_
rlabel metal1 17526 25942 17526 25942 0 _305_
rlabel metal2 17158 26282 17158 26282 0 _306_
rlabel metal2 15962 24718 15962 24718 0 _307_
rlabel metal2 15686 24412 15686 24412 0 _308_
rlabel metal1 16882 23800 16882 23800 0 _309_
rlabel metal1 16698 23664 16698 23664 0 _310_
rlabel metal2 17250 24854 17250 24854 0 _311_
rlabel metal1 17342 25840 17342 25840 0 _312_
rlabel metal1 17158 26010 17158 26010 0 _313_
rlabel metal2 18170 27778 18170 27778 0 _314_
rlabel via1 17618 28050 17618 28050 0 _315_
rlabel metal1 18262 28186 18262 28186 0 _316_
rlabel metal2 25438 34170 25438 34170 0 _317_
rlabel metal1 19228 34442 19228 34442 0 _318_
rlabel metal1 20056 35054 20056 35054 0 _319_
rlabel metal1 21252 34714 21252 34714 0 _320_
rlabel metal2 22034 34782 22034 34782 0 _321_
rlabel metal1 23138 34578 23138 34578 0 _322_
rlabel metal2 25254 34340 25254 34340 0 _323_
rlabel metal1 26404 34170 26404 34170 0 _324_
rlabel metal1 26818 34578 26818 34578 0 _325_
rlabel metal2 15870 19788 15870 19788 0 _326_
rlabel metal1 16606 22474 16606 22474 0 _327_
rlabel metal1 18584 21998 18584 21998 0 _328_
rlabel metal2 18814 22039 18814 22039 0 _329_
rlabel metal1 18446 21930 18446 21930 0 _330_
rlabel metal1 19550 26316 19550 26316 0 _331_
rlabel metal1 18722 23052 18722 23052 0 _332_
rlabel metal2 19826 27506 19826 27506 0 _333_
rlabel metal1 18814 27472 18814 27472 0 _334_
rlabel metal1 22218 27608 22218 27608 0 _335_
rlabel metal1 21160 26554 21160 26554 0 _336_
rlabel metal2 22402 28050 22402 28050 0 _337_
rlabel metal1 25070 16048 25070 16048 0 _338_
rlabel metal2 22126 15198 22126 15198 0 _339_
rlabel metal1 18032 14314 18032 14314 0 _340_
rlabel metal2 18354 14586 18354 14586 0 _341_
rlabel metal1 19136 14586 19136 14586 0 _342_
rlabel metal1 19918 14586 19918 14586 0 _343_
rlabel metal1 20286 14518 20286 14518 0 _344_
rlabel metal1 21850 14994 21850 14994 0 _345_
rlabel metal1 22908 15130 22908 15130 0 _346_
rlabel metal1 24978 16116 24978 16116 0 _347_
rlabel metal1 25392 16218 25392 16218 0 _348_
rlabel metal2 18722 33490 18722 33490 0 _349_
rlabel metal2 20838 33099 20838 33099 0 _350_
rlabel metal2 21298 33524 21298 33524 0 _351_
rlabel metal1 22908 33490 22908 33490 0 _352_
rlabel metal2 23322 33082 23322 33082 0 _353_
rlabel metal2 24058 33354 24058 33354 0 _354_
rlabel metal2 22402 32606 22402 32606 0 _355_
rlabel metal2 25070 31518 25070 31518 0 _356_
rlabel metal1 24610 31824 24610 31824 0 _357_
rlabel metal1 25530 31280 25530 31280 0 _358_
rlabel metal1 25254 31348 25254 31348 0 _359_
rlabel metal2 26818 32266 26818 32266 0 _360_
rlabel metal2 24564 45540 24564 45540 0 clk
rlabel metal1 20194 36074 20194 36074 0 clknet_0_clk
rlabel metal1 6394 16116 6394 16116 0 clknet_3_0__leaf_clk
rlabel metal1 4186 24786 4186 24786 0 clknet_3_1__leaf_clk
rlabel metal1 12236 13362 12236 13362 0 clknet_3_2__leaf_clk
rlabel metal1 24978 18122 24978 18122 0 clknet_3_3__leaf_clk
rlabel metal1 4646 29614 4646 29614 0 clknet_3_4__leaf_clk
rlabel metal1 9844 44914 9844 44914 0 clknet_3_5__leaf_clk
rlabel metal2 17802 34000 17802 34000 0 clknet_3_6__leaf_clk
rlabel metal1 19090 38794 19090 38794 0 clknet_3_7__leaf_clk
rlabel metal1 6072 29818 6072 29818 0 debounce0_a.button_hist\[0\]
rlabel metal1 7176 30770 7176 30770 0 debounce0_a.button_hist\[1\]
rlabel metal2 6762 30226 6762 30226 0 debounce0_a.button_hist\[2\]
rlabel metal1 7774 30124 7774 30124 0 debounce0_a.button_hist\[3\]
rlabel metal1 9338 29716 9338 29716 0 debounce0_a.button_hist\[4\]
rlabel metal1 10350 29274 10350 29274 0 debounce0_a.button_hist\[5\]
rlabel metal1 9062 30022 9062 30022 0 debounce0_a.button_hist\[6\]
rlabel metal2 10350 30294 10350 30294 0 debounce0_a.button_hist\[7\]
rlabel metal1 9982 25874 9982 25874 0 debounce0_a.debounced
rlabel metal2 5474 24412 5474 24412 0 debounce0_b.button_hist\[0\]
rlabel metal1 6348 24242 6348 24242 0 debounce0_b.button_hist\[1\]
rlabel metal2 7314 23358 7314 23358 0 debounce0_b.button_hist\[2\]
rlabel metal2 6394 24650 6394 24650 0 debounce0_b.button_hist\[3\]
rlabel metal2 6762 22848 6762 22848 0 debounce0_b.button_hist\[4\]
rlabel metal2 7038 19924 7038 19924 0 debounce0_b.button_hist\[5\]
rlabel metal2 6210 19652 6210 19652 0 debounce0_b.button_hist\[6\]
rlabel metal2 6854 21080 6854 21080 0 debounce0_b.button_hist\[7\]
rlabel metal1 8970 22644 8970 22644 0 debounce0_b.debounced
rlabel metal2 12190 44438 12190 44438 0 debounce1_a.button_hist\[0\]
rlabel metal1 12328 43826 12328 43826 0 debounce1_a.button_hist\[1\]
rlabel metal1 12006 44506 12006 44506 0 debounce1_a.button_hist\[2\]
rlabel metal2 12098 45220 12098 45220 0 debounce1_a.button_hist\[3\]
rlabel metal2 12466 43044 12466 43044 0 debounce1_a.button_hist\[4\]
rlabel metal1 14398 43418 14398 43418 0 debounce1_a.button_hist\[5\]
rlabel metal1 13938 44948 13938 44948 0 debounce1_a.button_hist\[6\]
rlabel metal1 13018 44506 13018 44506 0 debounce1_a.button_hist\[7\]
rlabel metal2 13478 39372 13478 39372 0 debounce1_a.debounced
rlabel metal1 8648 37434 8648 37434 0 debounce1_b.button_hist\[0\]
rlabel metal1 9384 36210 9384 36210 0 debounce1_b.button_hist\[1\]
rlabel metal1 10948 34714 10948 34714 0 debounce1_b.button_hist\[2\]
rlabel metal1 9384 36686 9384 36686 0 debounce1_b.button_hist\[3\]
rlabel metal2 9706 37536 9706 37536 0 debounce1_b.button_hist\[4\]
rlabel metal1 9200 39066 9200 39066 0 debounce1_b.button_hist\[5\]
rlabel metal1 10120 37910 10120 37910 0 debounce1_b.button_hist\[6\]
rlabel metal2 10626 38522 10626 38522 0 debounce1_b.button_hist\[7\]
rlabel metal2 12558 36924 12558 36924 0 debounce1_b.debounced
rlabel metal1 8050 9044 8050 9044 0 debounce2_a.button_hist\[0\]
rlabel metal1 10396 9418 10396 9418 0 debounce2_a.button_hist\[1\]
rlabel metal1 11086 11220 11086 11220 0 debounce2_a.button_hist\[2\]
rlabel metal2 10534 10285 10534 10285 0 debounce2_a.button_hist\[3\]
rlabel metal1 11086 10132 11086 10132 0 debounce2_a.button_hist\[4\]
rlabel metal2 9982 8500 9982 8500 0 debounce2_a.button_hist\[5\]
rlabel metal1 10396 9690 10396 9690 0 debounce2_a.button_hist\[6\]
rlabel metal1 11224 9894 11224 9894 0 debounce2_a.button_hist\[7\]
rlabel metal1 13754 14280 13754 14280 0 debounce2_a.debounced
rlabel metal1 5934 16558 5934 16558 0 debounce2_b.button_hist\[0\]
rlabel metal1 8694 16558 8694 16558 0 debounce2_b.button_hist\[1\]
rlabel metal2 8326 15742 8326 15742 0 debounce2_b.button_hist\[2\]
rlabel metal2 8510 15742 8510 15742 0 debounce2_b.button_hist\[3\]
rlabel metal1 10580 15130 10580 15130 0 debounce2_b.button_hist\[4\]
rlabel metal1 10166 16660 10166 16660 0 debounce2_b.button_hist\[5\]
rlabel metal1 9844 18054 9844 18054 0 debounce2_b.button_hist\[6\]
rlabel metal2 10350 15436 10350 15436 0 debounce2_b.button_hist\[7\]
rlabel metal1 12604 15674 12604 15674 0 debounce2_b.debounced
rlabel metal1 12185 20434 12185 20434 0 enc0\[0\]
rlabel metal1 12006 21930 12006 21930 0 enc0\[1\]
rlabel metal2 12374 25466 12374 25466 0 enc0\[2\]
rlabel metal1 14214 26996 14214 26996 0 enc0\[3\]
rlabel metal1 13892 32198 13892 32198 0 enc0\[4\]
rlabel metal1 14582 33388 14582 33388 0 enc0\[5\]
rlabel metal2 17526 33762 17526 33762 0 enc0\[6\]
rlabel metal1 16514 27370 16514 27370 0 enc0\[7\]
rlabel metal3 751 29308 751 29308 0 enc0_a
rlabel metal3 751 24548 751 24548 0 enc0_b
rlabel metal1 16882 39440 16882 39440 0 enc1\[0\]
rlabel metal1 18538 38828 18538 38828 0 enc1\[1\]
rlabel metal1 20838 40052 20838 40052 0 enc1\[2\]
rlabel metal1 21482 42738 21482 42738 0 enc1\[3\]
rlabel metal2 24058 39610 24058 39610 0 enc1\[4\]
rlabel metal1 24334 41446 24334 41446 0 enc1\[5\]
rlabel metal2 27738 40494 27738 40494 0 enc1\[6\]
rlabel metal1 27600 36550 27600 36550 0 enc1\[7\]
rlabel metal2 6578 48161 6578 48161 0 enc1_a
rlabel metal3 751 32708 751 32708 0 enc1_b
rlabel metal1 15134 11118 15134 11118 0 enc2\[0\]
rlabel metal1 15824 10778 15824 10778 0 enc2\[1\]
rlabel metal1 18906 10030 18906 10030 0 enc2\[2\]
rlabel metal2 20102 9214 20102 9214 0 enc2\[3\]
rlabel metal1 21344 14314 21344 14314 0 enc2\[4\]
rlabel metal1 23276 12818 23276 12818 0 enc2\[5\]
rlabel metal2 25990 9588 25990 9588 0 enc2\[6\]
rlabel metal1 25944 13498 25944 13498 0 enc2\[7\]
rlabel metal2 5198 1027 5198 1027 0 enc2_a
rlabel metal3 751 15708 751 15708 0 enc2_b
rlabel metal1 10212 23766 10212 23766 0 encoder0.old_a
rlabel metal1 10396 23290 10396 23290 0 encoder0.old_b
rlabel metal2 14582 39100 14582 39100 0 encoder1.old_a
rlabel metal2 14306 37468 14306 37468 0 encoder1.old_b
rlabel metal1 13570 14348 13570 14348 0 encoder2.old_a
rlabel metal1 13938 15062 13938 15062 0 encoder2.old_b
rlabel metal1 3082 29648 3082 29648 0 net1
rlabel metal2 28290 16252 28290 16252 0 net10
rlabel metal1 23230 17204 23230 17204 0 net100
rlabel metal1 23000 32402 23000 32402 0 net101
rlabel metal1 19504 23154 19504 23154 0 net102
rlabel metal2 21574 27676 21574 27676 0 net103
rlabel metal2 24978 31484 24978 31484 0 net104
rlabel metal1 24932 31790 24932 31790 0 net105
rlabel metal2 25622 17408 25622 17408 0 net106
rlabel metal1 26726 32912 26726 32912 0 net107
rlabel metal1 16560 22610 16560 22610 0 net108
rlabel metal1 19136 16558 19136 16558 0 net109
rlabel metal1 28014 23290 28014 23290 0 net11
rlabel metal2 19090 27268 19090 27268 0 net110
rlabel metal1 27646 37230 27646 37230 0 net111
rlabel metal1 17710 22678 17710 22678 0 net112
rlabel metal1 21206 32810 21206 32810 0 net113
rlabel metal2 18170 15776 18170 15776 0 net114
rlabel metal1 17756 15674 17756 15674 0 net115
rlabel metal1 24702 13260 24702 13260 0 net116
rlabel metal1 23000 17646 23000 17646 0 net117
rlabel metal2 20378 35190 20378 35190 0 net118
rlabel metal1 20102 17612 20102 17612 0 net119
rlabel metal1 24794 12750 24794 12750 0 net12
rlabel metal1 22126 27540 22126 27540 0 net120
rlabel metal1 13570 32878 13570 32878 0 net121
rlabel metal1 16054 19380 16054 19380 0 net122
rlabel metal1 19090 33082 19090 33082 0 net123
rlabel metal1 19964 32538 19964 32538 0 net124
rlabel metal2 20838 42058 20838 42058 0 net125
rlabel metal1 19918 9044 19918 9044 0 net13
rlabel metal1 20286 38386 20286 38386 0 net14
rlabel metal2 21206 39916 21206 39916 0 net15
rlabel metal1 13708 32402 13708 32402 0 net16
rlabel metal2 11914 32096 11914 32096 0 net17
rlabel metal2 17250 33184 17250 33184 0 net18
rlabel metal1 12098 22202 12098 22202 0 net19
rlabel metal1 2714 24718 2714 24718 0 net2
rlabel metal1 10212 17646 10212 17646 0 net20
rlabel metal1 6072 15470 6072 15470 0 net21
rlabel metal1 3588 24174 3588 24174 0 net22
rlabel metal1 9348 18258 9348 18258 0 net23
rlabel metal1 6578 35734 6578 35734 0 net24
rlabel metal1 13800 43758 13800 43758 0 net25
rlabel metal2 8326 39865 8326 39865 0 net26
rlabel metal1 12650 37774 12650 37774 0 net27
rlabel metal1 18676 16150 18676 16150 0 net28
rlabel metal2 22126 18156 22126 18156 0 net29
rlabel metal1 6946 47158 6946 47158 0 net3
rlabel metal1 23690 18734 23690 18734 0 net30
rlabel metal2 20194 41344 20194 41344 0 net31
rlabel metal2 20930 33490 20930 33490 0 net32
rlabel metal1 26588 41582 26588 41582 0 net33
rlabel via2 28566 19805 28566 19805 0 net34
rlabel metal2 27094 1588 27094 1588 0 net35
rlabel via2 28566 27931 28566 27931 0 net36
rlabel metal3 751 30668 751 30668 0 net37
rlabel metal3 751 28628 751 28628 0 net38
rlabel metal3 751 31348 751 31348 0 net39
rlabel metal1 2576 33082 2576 33082 0 net4
rlabel metal3 820 9588 820 9588 0 net40
rlabel metal2 28198 15793 28198 15793 0 net41
rlabel metal3 751 32028 751 32028 0 net42
rlabel via2 28566 22525 28566 22525 0 net43
rlabel metal1 12696 42534 12696 42534 0 net44
rlabel metal1 12507 40018 12507 40018 0 net45
rlabel metal1 11500 16490 11500 16490 0 net46
rlabel metal1 10902 29478 10902 29478 0 net47
rlabel metal2 11730 11764 11730 11764 0 net48
rlabel metal2 12926 10914 12926 10914 0 net49
rlabel metal2 5474 5542 5474 5542 0 net5
rlabel metal2 10810 17170 10810 17170 0 net50
rlabel metal2 11086 16082 11086 16082 0 net51
rlabel metal1 11224 36822 11224 36822 0 net52
rlabel metal2 10166 37808 10166 37808 0 net53
rlabel metal2 10534 37230 10534 37230 0 net54
rlabel metal2 11914 44268 11914 44268 0 net55
rlabel metal1 11776 8942 11776 8942 0 net56
rlabel metal1 7314 21114 7314 21114 0 net57
rlabel metal2 8142 22882 8142 22882 0 net58
rlabel metal2 6486 31076 6486 31076 0 net59
rlabel metal2 3266 15674 3266 15674 0 net6
rlabel metal2 11822 43724 11822 43724 0 net60
rlabel metal2 9430 9316 9430 9316 0 net61
rlabel metal2 8142 24650 8142 24650 0 net62
rlabel metal1 10120 38386 10120 38386 0 net63
rlabel metal2 8510 39610 8510 39610 0 net64
rlabel metal2 7222 23868 7222 23868 0 net65
rlabel metal2 8602 38148 8602 38148 0 net66
rlabel metal1 9568 10574 9568 10574 0 net67
rlabel metal1 9844 14450 9844 14450 0 net68
rlabel metal1 8096 14382 8096 14382 0 net69
rlabel metal2 28382 9282 28382 9282 0 net7
rlabel metal1 8510 29172 8510 29172 0 net70
rlabel metal1 5520 30770 5520 30770 0 net71
rlabel metal2 8786 18700 8786 18700 0 net72
rlabel metal2 11362 11084 11362 11084 0 net73
rlabel metal2 7314 29580 7314 29580 0 net74
rlabel metal1 5704 29274 5704 29274 0 net75
rlabel metal1 8556 31246 8556 31246 0 net76
rlabel metal1 15088 44914 15088 44914 0 net77
rlabel metal1 8648 36686 8648 36686 0 net78
rlabel metal2 7590 8636 7590 8636 0 net79
rlabel metal1 28336 31790 28336 31790 0 net8
rlabel metal1 6256 20434 6256 20434 0 net80
rlabel metal2 6946 19482 6946 19482 0 net81
rlabel metal2 8970 35836 8970 35836 0 net82
rlabel metal2 6026 23868 6026 23868 0 net83
rlabel metal1 14030 43758 14030 43758 0 net84
rlabel metal1 8924 44302 8924 44302 0 net85
rlabel metal2 11178 8908 11178 8908 0 net86
rlabel metal1 4692 24242 4692 24242 0 net87
rlabel metal2 6302 15980 6302 15980 0 net88
rlabel metal2 5842 16252 5842 16252 0 net89
rlabel metal2 28290 35462 28290 35462 0 net9
rlabel metal1 8326 44404 8326 44404 0 net90
rlabel metal2 6394 35428 6394 35428 0 net91
rlabel metal1 17986 34000 17986 34000 0 net92
rlabel metal1 17388 17170 17388 17170 0 net93
rlabel metal1 15594 18258 15594 18258 0 net94
rlabel metal2 21022 17340 21022 17340 0 net95
rlabel metal1 25760 17714 25760 17714 0 net96
rlabel metal1 26986 16490 26986 16490 0 net97
rlabel metal1 26450 34578 26450 34578 0 net98
rlabel metal1 27411 35054 27411 35054 0 net99
rlabel metal2 16146 19431 16146 19431 0 pwm0.count\[0\]
rlabel metal1 16238 20434 16238 20434 0 pwm0.count\[1\]
rlabel metal1 16330 21862 16330 21862 0 pwm0.count\[2\]
rlabel metal1 18906 22066 18906 22066 0 pwm0.count\[3\]
rlabel via1 16879 25874 16879 25874 0 pwm0.count\[4\]
rlabel metal2 17986 27948 17986 27948 0 pwm0.count\[5\]
rlabel metal2 19458 28390 19458 28390 0 pwm0.count\[6\]
rlabel metal1 16882 27574 16882 27574 0 pwm0.count\[7\]
rlabel metal3 28896 31348 28896 31348 0 pwm0_out
rlabel metal2 18630 35156 18630 35156 0 pwm1.count\[0\]
rlabel metal1 18722 33830 18722 33830 0 pwm1.count\[1\]
rlabel metal1 19596 33286 19596 33286 0 pwm1.count\[2\]
rlabel metal1 21482 34544 21482 34544 0 pwm1.count\[3\]
rlabel metal2 22954 34170 22954 34170 0 pwm1.count\[4\]
rlabel metal1 24311 34578 24311 34578 0 pwm1.count\[5\]
rlabel metal2 25622 34238 25622 34238 0 pwm1.count\[6\]
rlabel metal2 28014 34272 28014 34272 0 pwm1.count\[7\]
rlabel via2 28474 35445 28474 35445 0 pwm1_out
rlabel metal2 18262 14960 18262 14960 0 pwm2.count\[0\]
rlabel metal1 17434 14994 17434 14994 0 pwm2.count\[1\]
rlabel metal1 19734 17068 19734 17068 0 pwm2.count\[2\]
rlabel viali 20380 15470 20380 15470 0 pwm2.count\[3\]
rlabel metal1 21160 15470 21160 15470 0 pwm2.count\[4\]
rlabel metal1 23552 18394 23552 18394 0 pwm2.count\[5\]
rlabel metal1 24288 17578 24288 17578 0 pwm2.count\[6\]
rlabel metal1 26450 18054 26450 18054 0 pwm2.count\[7\]
rlabel metal2 28474 16303 28474 16303 0 pwm2_out
rlabel metal2 28566 8347 28566 8347 0 reset
rlabel metal2 28474 23341 28474 23341 0 sync
<< properties >>
string FIXED_BBOX 0 0 30000 50000
<< end >>
