VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rgb_mixer
  CLASS BLOCK ;
  FOREIGN rgb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 246.000 122.730 250.000 ;
    END
  END clk
  PIN enc0_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END enc0_a
  PIN enc0_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END enc0_b
  PIN enc1_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 246.000 32.570 250.000 ;
    END
  END enc1_a
  PIN enc1_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END enc1_b
  PIN enc2_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END enc2_a
  PIN enc2_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END enc2_b
  PIN io_oeb_high[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 112.240 150.000 112.840 ;
    END
  END io_oeb_high[0]
  PIN io_oeb_high[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 98.640 150.000 99.240 ;
    END
  END io_oeb_high[1]
  PIN io_oeb_high[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END io_oeb_high[2]
  PIN io_oeb_high[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 139.440 150.000 140.040 ;
    END
  END io_oeb_high[3]
  PIN io_oeb_high[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END io_oeb_high[4]
  PIN io_oeb_high[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END io_oeb_high[5]
  PIN io_oeb_low[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END io_oeb_low[0]
  PIN io_oeb_low[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END io_oeb_low[1]
  PIN io_oeb_low[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 78.240 150.000 78.840 ;
    END
  END io_oeb_low[2]
  PIN io_oeb_low[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_oeb_low[3]
  PIN pwm0_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 156.440 150.000 157.040 ;
    END
  END pwm0_out
  PIN pwm1_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 176.840 150.000 177.440 ;
    END
  END pwm1_out
  PIN pwm2_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 81.640 150.000 82.240 ;
    END
  END pwm2_out
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 40.840 150.000 41.440 ;
    END
  END reset
  PIN sync
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 115.640 150.000 116.240 ;
    END
  END sync
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 236.880 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.760 144.630 236.830 ;
      LAYER li1 ;
        RECT 5.520 10.795 144.440 236.725 ;
      LAYER met1 ;
        RECT 4.210 10.640 144.440 236.880 ;
      LAYER met2 ;
        RECT 4.230 245.720 32.010 246.570 ;
        RECT 32.850 245.720 122.170 246.570 ;
        RECT 123.010 245.720 142.970 246.570 ;
        RECT 4.230 4.280 142.970 245.720 ;
        RECT 4.230 4.000 25.570 4.280 ;
        RECT 26.410 4.000 135.050 4.280 ;
        RECT 135.890 4.000 142.970 4.280 ;
      LAYER met3 ;
        RECT 3.990 177.840 146.000 236.805 ;
        RECT 3.990 176.440 145.600 177.840 ;
        RECT 3.990 164.240 146.000 176.440 ;
        RECT 4.400 162.840 146.000 164.240 ;
        RECT 3.990 160.840 146.000 162.840 ;
        RECT 4.400 159.440 146.000 160.840 ;
        RECT 3.990 157.440 146.000 159.440 ;
        RECT 4.400 156.040 145.600 157.440 ;
        RECT 3.990 154.040 146.000 156.040 ;
        RECT 4.400 152.640 146.000 154.040 ;
        RECT 3.990 147.240 146.000 152.640 ;
        RECT 4.400 145.840 146.000 147.240 ;
        RECT 3.990 143.840 146.000 145.840 ;
        RECT 4.400 142.440 146.000 143.840 ;
        RECT 3.990 140.440 146.000 142.440 ;
        RECT 3.990 139.040 145.600 140.440 ;
        RECT 3.990 123.440 146.000 139.040 ;
        RECT 4.400 122.040 146.000 123.440 ;
        RECT 3.990 116.640 146.000 122.040 ;
        RECT 3.990 115.240 145.600 116.640 ;
        RECT 3.990 113.240 146.000 115.240 ;
        RECT 3.990 111.840 145.600 113.240 ;
        RECT 3.990 99.640 146.000 111.840 ;
        RECT 3.990 98.240 145.600 99.640 ;
        RECT 3.990 82.640 146.000 98.240 ;
        RECT 3.990 81.240 145.600 82.640 ;
        RECT 3.990 79.240 146.000 81.240 ;
        RECT 4.400 77.840 145.600 79.240 ;
        RECT 3.990 48.640 146.000 77.840 ;
        RECT 4.400 47.240 146.000 48.640 ;
        RECT 3.990 41.840 146.000 47.240 ;
        RECT 3.990 40.440 145.600 41.840 ;
        RECT 3.990 10.715 146.000 40.440 ;
  END
END rgb_mixer
END LIBRARY

