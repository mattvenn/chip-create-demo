VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rgb_mixer
  CLASS BLOCK ;
  FOREIGN rgb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END clk
  PIN enc0_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 25.850 246.000 26.130 250.000 ;
    END
  END enc0_a
  PIN enc0_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END enc0_b
  PIN enc1_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END enc1_a
  PIN enc1_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END enc1_b
  PIN enc2_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END enc2_a
  PIN enc2_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END enc2_b
  PIN io_oeb_high[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 156.440 150.000 157.040 ;
    END
  END io_oeb_high[0]
  PIN io_oeb_high[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 136.040 150.000 136.640 ;
    END
  END io_oeb_high[1]
  PIN io_oeb_high[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_oeb_high[2]
  PIN io_oeb_high[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 246.000 122.730 250.000 ;
    END
  END io_oeb_high[3]
  PIN io_oeb_high[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_oeb_high[4]
  PIN io_oeb_high[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END io_oeb_high[5]
  PIN io_oeb_low[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_oeb_low[0]
  PIN io_oeb_low[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_oeb_low[1]
  PIN io_oeb_low[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 71.440 150.000 72.040 ;
    END
  END io_oeb_low[2]
  PIN io_oeb_low[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_oeb_low[3]
  PIN pwm0_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 246.000 109.850 250.000 ;
    END
  END pwm0_out
  PIN pwm1_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 159.840 150.000 160.440 ;
    END
  END pwm1_out
  PIN pwm2_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 78.240 150.000 78.840 ;
    END
  END pwm2_out
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 146.000 40.840 150.000 41.440 ;
    END
  END reset
  PIN sync
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 85.040 150.000 85.640 ;
    END
  END sync
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 236.880 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.760 144.630 236.830 ;
      LAYER li1 ;
        RECT 5.520 10.795 144.440 236.725 ;
      LAYER met1 ;
        RECT 0.530 10.640 144.440 236.880 ;
      LAYER met2 ;
        RECT 0.550 245.720 25.570 246.570 ;
        RECT 26.410 245.720 109.290 246.570 ;
        RECT 110.130 245.720 122.170 246.570 ;
        RECT 123.010 245.720 142.510 246.570 ;
        RECT 0.550 4.280 142.510 245.720 ;
        RECT 0.550 4.000 28.790 4.280 ;
        RECT 29.630 4.000 109.290 4.280 ;
        RECT 110.130 4.000 142.510 4.280 ;
      LAYER met3 ;
        RECT 0.525 222.040 146.000 236.805 ;
        RECT 4.400 220.640 146.000 222.040 ;
        RECT 0.525 191.440 146.000 220.640 ;
        RECT 4.400 190.040 146.000 191.440 ;
        RECT 0.525 160.840 146.000 190.040 ;
        RECT 4.400 159.440 145.600 160.840 ;
        RECT 0.525 157.440 146.000 159.440 ;
        RECT 0.525 156.040 145.600 157.440 ;
        RECT 0.525 150.640 146.000 156.040 ;
        RECT 4.400 149.240 146.000 150.640 ;
        RECT 0.525 147.240 146.000 149.240 ;
        RECT 4.400 145.840 146.000 147.240 ;
        RECT 0.525 137.040 146.000 145.840 ;
        RECT 0.525 135.640 145.600 137.040 ;
        RECT 0.525 120.040 146.000 135.640 ;
        RECT 4.400 118.640 146.000 120.040 ;
        RECT 0.525 116.640 146.000 118.640 ;
        RECT 4.400 115.240 146.000 116.640 ;
        RECT 0.525 109.840 146.000 115.240 ;
        RECT 4.400 108.440 146.000 109.840 ;
        RECT 0.525 89.440 146.000 108.440 ;
        RECT 4.400 88.040 146.000 89.440 ;
        RECT 0.525 86.040 146.000 88.040 ;
        RECT 4.400 84.640 145.600 86.040 ;
        RECT 0.525 79.240 146.000 84.640 ;
        RECT 0.525 77.840 145.600 79.240 ;
        RECT 0.525 72.440 146.000 77.840 ;
        RECT 0.525 71.040 145.600 72.440 ;
        RECT 0.525 41.840 146.000 71.040 ;
        RECT 0.525 40.440 145.600 41.840 ;
        RECT 0.525 10.715 146.000 40.440 ;
  END
END rgb_mixer
END LIBRARY

